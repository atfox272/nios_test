// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
JweQU8k2648wuj38P4MLnD5Bh0MQclxMdUc+AgKKTHovYqlnvf39c+Wm8CFNeRy6QfonScE5I7SI
jVZuJNJ6FiAjR3lNbpsAejvdFth7sJf/XJLIS1ur0SWFddBxtwcMAux+sFUa1HhdCCCvkB9gAahQ
Y6FpztuW1+Y/plZ2//ACYn94fALpLjWx7bxkxmUdMc7eGlxd2YEnYVWdTi5fr2q0DaVnmrTIqXIn
wsf8jQB6/aiAWAobTRS06oHOCrG5iZCTaBUhxQB31QsNDrGZT4rUEUrR6zoKnWuGVFCNRx8mrjul
UzIxnwc0SDMPe1SxH0NZSlaVVPj8NSSRNF8Jog==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6272)
lObkLcxVAZmmtsv8LuhzkNPcylFyep5MLTPVP3mV014D8R9RZRhICX8zUEOpiqHLGtjX1G588GLb
DMCsIiuEhxOhMfXVfz9w9XpVc2Vy1EkK3WuyRIec8FIqwDF1cxxxQR6QHIc5v2L8ZMqyIMc7UgJq
tLZXij9DlDS3bctzGc6nyvCX+gZZtDRmQQJC9NFC0DLzd11aX2M6q5ZZbUPegiBty8tZDTwHWER/
2qXjKA+Aps+iamI5J3NizzxEZUi96U1NrIFSqrI33EAqhMBREJ8Q7c3jlE0qVHZFswuH0FotYqy3
rwiz0nT+lw9VXx7cCl0Of4F6TOHhpKxD9afksOjymyYM5pIccZ/UmPbLj5hIJNCmJJDMttf4Hmzv
Y0sD65Vm0orcVShlld9iVequBc/znFTfuAUKJeLQxjKdVCEY/Pvqyf4TjiXLYQnI5Zq72kMH+TEx
+xLW4dra/tiBSLQav6CnamEXMarD97csa4mbLdVi+/rTJJpQRXQ18Is32XVS2AaiwtII6bxUpA+0
ygLvB1APHk/U0uFY/OBeYFwd7TY/YROx5pA0whRtFa6h5sLBZn5sKLsw4m5852zQeqXb/Qfn7kXB
fCocSGAMxowMV9npUHWBusSYQRp6/5JxW3F/r720th0/9Bc0WC731IbijlLF3q9AUrtIZ7jndkT6
ZpC4PLgFjephHq1qr2WG+p+/zGaYOns+JH2yqjXI/6uY8ho+Jym5PP9kq1Omwtl3gmHWaDqAdokQ
4NU2y3PTqtUl3l7Rqc1CjIFfw2x1/2gJlag7Dr/zpdnrTBNdPS6UGhvNpoGJ1SQZnTT1ZhxfFO69
gsvIqvIVpq9N0opDHMKCuRhDVLP0hpdQ8eRRy3bob9rrDZOy11jboTYM6tVoKL2IY5cjMi/z6rIy
TFjXT+QiFztWxKRjueVxEr0Xe/gNVQ34voWTYWncKsvRUA1p3f5YQeJ/iVLY8J/4tbEbZjzIXUPs
4UWF3ynwC7GtXJqO07JEhCyjE9cR3Zq+ee8MAMlrhzcWW1hsHpvpsjbcCHMZMKnYvn+5yi9O7DhQ
pA7uIiKeOE8x0kj9jAL2WxaCGeTwYlJB4CWzAxXsO0OnuawN8XyyymWdNVINg50PhjM8pV8BTOA1
uH3BrKWowHYyscAbo2cnp51BF8Pb9EDo9LGmRf6NBy1w/Uzgf5OITjSeZ7Pr/hAylre2qB2Zjjhj
ZRNvnR8nEEPA2AeqlIZKwsa0QuUjwPclq6Cuhx/iVduSQJZH5UaCFQoLcUjAiIVBBzLJk2Kf9df9
tBnLDXnhC4sBK2oyh+0XM/10bXc3tTA+x8GB3L5lUcbuPb5DFMcgPobG/QJZ/os/KtTYF6b2VslX
rERRCwPlu0uyhJGnPCG5bLKOHKIZmLCJ2LQanN8C8adK+bX6Yv0REa1g3wyuu7G9LfvtknhtkaSf
nkoyi8avqBYcxzecuj6mAPD8pdTEzt1BnrQ8xSmF/08Z/zdG78c7ZaF+Emhbt/LiihNRV0+QiNZX
lcwhB/rn7W0U62PDdbgHGTmMIQEvBeIDHkaWaVzrjJ+Ci+p9q0eGSCfictcQ6Jdl6m6zmWpHmPu3
swC2dCP5GngwBrOq2ZTEdfx4gKUY0ECGYRySfwYjv40+9H3xgEkbdwbjnKE7uYMSTLs8EYWPA7jU
obkAVrDCpYbk4hkNfpFRtLo8QwJPoJorgN2bXy5GtwpGSTxfqBM22KYvtX9pPHOyMZ2FSdhIV+ac
tZaQ2oYE3wnU1CxxYzhe7vLPowyIdyE/QaxPRF7VJQ/FDKU5ZoyVvptySA+CY/V2G1i9rPc1icI9
vJewoVXzeDnfRNEwBFzpM6DObCt//eNEAC7uC0VbMqk9e5HEEW+vN/64vJ6efOgrnspeODd1/vuH
/l/TA2dpbUFMNlb75GJqLoSa16nL3r2F/oyzGULUlHtHIy/Ex4W0nVa96DapSutElGrVlW81xQ3a
uAmdi4tauzUGrtF4DEfUPdjTlLMzNqQ3UHvWo0ILbcFdwA04sPMA9sH0oyE/Mjgi/5NjFXIsJUk7
jAxYPgGoFKZSXZebn/JcrCZQFiG+q4PlBu8C8JrAolSQHDCC1OO+KU8/PgZJocwKTJE6ZrjBxWyP
aVKBmpCjEaMdg49hbh0DK/HMXEwmtWh41mUQVZr2gcm9sY/hHy8v61SkjTmUX9gf22qtBuH19TVw
m3zGGJvyMqkEszS8USgFFMn6Dps86fk/iAAH9cRhe4IE3XIA0Ai3H4Fes5siSAkY8alMXC775QdK
BZo74s6mAYywIjqEbw6gfcySidhWRj38X3tWNica5X28tPyv47moCnEPCibt339BUv+UZAwtoIuh
hFYdbblRmcC9trfkDTeJwrVrkNSB5dswvotitt4MszEO5XUdUr/NITSlIbb6jCqGLOAb0c0tN6nA
ZOGvwQS3KsYgfl+4HueK9iZdWXN9pcoO+KpkbwT4aG/f7icSnUVwrnM+vVYqlt1whS8/UQT5kVNw
hyn5KG+n4f+MYSqsooBSAGZO3muziBbHnXa2p65gMAQKwoPFZ3PN9xwVJ+KGMf8Vtp+V2GKSMs3I
j4h5/u9FT24ZddkqUHo0K8W8MIR3loQg2JV10nuCGpfGP5c15iMQ7hFgGWE3ygPFg5c/BGjncZZv
+u4HYbTdFQXJg6HN6XnDC8UN/Q+KKwWdrxjjx0IOhVjgSrvvJMYItTrfjSUnf2pna2fH5ewDUvmG
iNpWJFhffLMPo/XuSIXD+h9vcLnv/1Ak2N8X8a9jWE5rzDU6ZL7W8gZkOdJVmXtgw1J7l+KpTeGb
1eJR2q/XiyZWwD2wgpvIVMd/J2UAKgDIYUG77Rfkc28GlPgJ1+DTgw/ovLDuIefD/IlY5wLtLzZu
Yv6OuB9Ji6LZlzCHhAFRC0ftGiP5cLnubULjP1n9mHVEICyATBTW31n+97W5DQqfZQVejlrVN+zq
O437SwClcdbRVHCULETQNT9RF043SmsEMNYQ4/pltRswaW5H82i3SAHzIAxUSmHoYdENpUkA3qfk
D7l+s6wNZywj9T0/fiEfLe9GG7AVzeHboOp+znIO6AJ8rHtKH8C0YNd4PmulfkoZizjbzfPeDAFQ
Bsv0pJ9mnKARZAMAPzV48H0Xoh/12Sg+FsB6jung6iKBzfGxOPIajysoQlQILM+oSPYnQzHc/8/M
xjYQvv+5GAd7dL1K3wiZNq3JhEXi2clnDN51h91Z5qeN/UqlnfkXabA6NcJLKXb/HHgesFV1ID74
ZU9zognCCHVpYEz8C5p9IBFoIs7zAQurjsrYhPP3J1ITA0+KC6h/AMrfE8dOtyAZGtn4XiZ5XfV6
5VGhcl2KJfdM2JxPqNl00Q+23kDPQlDHaqWGZP7hcckK5VPM8OKh2inNwJB3tq3wvcjDiybXjoUt
vlTl3rqgUENVnunSBhkQsDQOjZ6L7Nt6lf2MGNZRKQGyouI71X5T18Lq4W2ioXKfWn5URXRcsjhd
qwRhETy4+BGP43UBnENwKLjMKilP07PCfsEll68ylKwq+uaeQLMf97zJ02HeQ0AS2bk0hhQVoPYB
tB1+hVH56HUt1HRnl0Et3chUNf1pgFft24NBbZwtBi5wxlzuGz4rs8er9FEIsLIHx2vo/kTAzTNm
8Nj2XKm6C95VJlW8T6tvLD1KXkIZzfhQ1dwwb9NfQMFKfnyHN7EMBWAyVeDD7cCxhQeiLuGzexlE
tyAVS+Srndk9Po/4pyXe0AxWjio5LGLWEkmyOddaerPnWPvj8eNvyEclOfQuKFxJ4VdT1hv0ioBH
plyYR80rfwm/8Oo7YH1X6nbynkXLwI+tgES9mRG3gvbdUrQOgL2D3d0e7gtA+iv5YyZXqgC/4qWk
heIdyg63s3nVNXmLSoKjHeMW9ObJ0Dy8i49OIgYf4NduncFBRLsPupG+wPnMgc41DcMKDJ67Q/zP
O5sfeP4urdNn+rHgGmTLZw8HtPNWce733HTSYoxcJJdo6WBMHLQh1QD/Y4GAPNZvlW/cmS/Jo5mW
kldP/YyqKVA6bdzTeJ2WOFapTUWnmxnQ6V2AD0gvAvc3cL1vYfElrrRo7nuabguotpzX7b44FpYg
LZLlTqyyB6TaGtVxFpAa2+GaQ4lhOsGJ9fghF8rOEWOQZFGPtDBUCZEiHSzTWyGqqdCVa2K7G77g
XF8aH6ohKrqKqFDjd6WZhbt0NyONZqMKcQ7OuGwVk3bIiVvPYdqYKCd6eoqdzyRtSC6baIcKaYvw
Jh6f3F99BU6Ff4sKdrywEGB7ByM18sS28RjVGqCyvo5ReXVuRoxysGUyy9K8tjuyAXC11/DLzBUQ
CBuuNOI1YQR6/HvTpIPrXaVGuCy0IMVlCJgbVHbCp1Q0Xd6J0eD6Pg/C1eFfo9J1SX7GogZenIzB
k/rI+Jks/oRzdzHr/2wXK7l6ihTBS9SGqSzZYRchCqsv6wfWL5noNadCWNC/UkYU+sm5roHx9W65
vis9pyjXLSSGB3JhR7AWsfZ+CbPlfKsU79NisSwVELBezKoA2Ab/eksb9cTGpoY4dRSLILl8veyG
eLi9dsXtQACheAFbbzHvxC7BK9q+2+DuMVgX8xaZP7wkrL99G5dWKij1LkKzy/Raa2ypmdf9pnUp
055XRfszD04BHtnXhopSNv2KFXovA51x8NClcm9PzwxdI44mcdClxQgyzCBOJPJyfi755u6KZTlx
9pO7R1JxduAy6z7Cd3sgigQPpMNp8f7HvtLjZ6QFMSaNc/gTqiDp1qhnJ56u2lh85heFYuehcY8w
XCCoJnLKyDujjZjFUz7QM+OsPCOBXJ7kR3+y4X6qay7YTMbxQPhnhkXbWZ20eW49115EG4ihlfEf
uXic0RRqKiceXPV29LVgbLJQxY8Ka8m3TBK8ZvKnt8TaoZzt/EJ1evFHKCazXTPzynxW44+saJ/b
B0PJF+EvejdgqjL3kvFh3+7PrAkX/GF6tJeHOFU4PgpPwQ6ISCWkFK/GB31SoXSF7fCoYi9aYkaB
9g0qH+bEW11wa/2c9Qc6nLc6CdIdjK9ktlf1xnVZurflkJ1Irxl6j+3bKCS5O0v6VVKQbia29y6z
89QzrKGDGP1ZDC0XI6nTTMaiRt3thYkgFMNjH1HOh8ulRDzA9g+9l/is0WwQziHPPyOyg0ENNjNy
JEE3eNTpxh8XwEwpefXbmRocXJkSKwjos7Zvq7fyNi0jjapGrR6rDWbvW+L6ucpLBBiulTq3ati/
Xb4/i1qDKDfmtcljCE/Mlm8OVaXMj2ZSO09bufAMA73QVfvL/YwoiiL0lJhcQnEj70nP5BkOFa56
JK8v+DSglAd6/BCwnxzb6bNhqikg3QLdV4rjhOurOwrJ+Q8R/0fysjmJFD2PRpRCoctKUnBX/URP
3SBqhW6CoXdTMGVeSIBpnmYlfqxR2YzoC27lTh+EvXlEZXE9zkncKq+YAOjbh5yJa8Jd/SJti4Yf
ggjXbTTL6wynTMU5uwWFm7m+yR4JFvIpMhVabBWOu0gqVyHeP5A+J04FKbYNntuxfEnXECA1AS1O
kOoEOAK3KZkNsR2uJzgr6Cuo6yrdM8AyML2FtAcXQEtTWiFxL9QDodbkfBYfcOmdXTI1TIELTzkj
lmm5h/SMD59zcVocV5jwG7uZVQjC9gJjjJDucKoBCl1JWPoSxauuLrexwrt5clLUFM88O1CbIZPN
KXxnduu4wfJ4xmjDQDnPZ7Bc6F9ZwgJtLBzbk8Bv0hG+u5wazFAN11ruyBdfG26hDTTQQyH9uAIK
IAgMd0cBVtGFBHVbyx9NhJjf8qgJl2Yy7kfpLVDPcQVB3MZ3alXEG9IanCSsi1mCDnYHqWQnWGUe
6caeWXyzn0DUP3vdDf36qbIvvFx7LcjgCxuqXXi8TUiYHbSmsVKvGwrKMJuifPBJ/y7IPd1A2Hhg
NuwdWoZ2mYPkxyL+72yokSeXt4Tg+2Z1FakBCaIY5AD6Vo//OI+QIcJreAfbxQKdmOU421CVAwnR
ZWLPbCjWmhA/UsRyiM0bP9CTNajLFkKY/P6SUBvZJ1RzXK/Zi32dFbWaULWjx9a9Mq2Jull47lkl
sgccgXh+Dp4z0Xgwty36KaBBPIp/uwuouY3nl3lbB2WfytmDc2dJnkzrC+igWRPJ80Why1N61XHW
hcW52Kh7D+1kgKM4imrq5S0i7mVbjFYDxd3kuqM/2fqizC9R1tjR1TdANZKRP0mUaIDP4yHayhFw
uehyUXsmZIuCPPJoX/AyusW426QmbelPAzU0OzkYpkaNU7GKVOlO1q6cwFwfi2yZQbNK8MkjwPwJ
izekCkJDCr0GUfKqmzesSsQeSmceCGK6exnOjU5VqCux7cKu11nC0D9TMQ+1bOziBfPhldADZeyV
4dCBPaJ/SkGBXv+MZzbLSHSq8OmplTPwhAIVfaDI8CBXru9AErG4NGlb2GuQZrdKOzVfUGa6wf+k
h8QJtI1DSqGeo6xo5LAyEaj7eQASiXY7zXju8QwI2qmrqV7MSxIWjdcYAKd6VEpG5SuWLYnYMhQw
X6HmfC+mheRZANOfGtkctx1Z3wkGtSTAptYqlFNs+52PyW+2UCqbxgi8VVyX++rrWMhLw5SBiZqF
gnc2htS+OZRVv4azYj93iwEzx2fUvopfu60KE/Zl8R+5XfOKPySPfxDq4qU1TfjZsnBVwLbWCl5Z
HD33j1ufTrqmmMgYaDWqTE3g3Ipi+OakyuW7XXkoiDfPkljIqjUSLlAhPLYButS2Jb3WPEQYw+1A
qS5XRTi8932zXhG0OP4XUXdGkdC3yGyT0Qh43PlO+5ULlR/iOrTiHy/wrJ92Jzk8A6QhekyYhRoB
aem5B6SqRKf9bGJENb8nToR18qJxEHM3pPxjDYzsJ1aBB/xvZ/MJcJb3yKksETGZ/3EswzgGZlMp
tf7/LhuXZX6ztH5YTbg5wahnTnCP4FgtpyujhmCBPEgYcxUiDPronFS+5YrUFlESiUQjfmBluWY9
xukB3p91yEhyy0Y1wr4Ql4Xh/TgqkAHCzTvvOTW5qai0s4/afA/isWdJFTY0S1Ttf9kaPbil51i3
BH3Ea6AHOTh3e00wpcEg/gCGnEkce5uFPbJgVN/UtZ3D8dNyZjLx86qS38PZpVKTqdWhAidgo8MK
d8yuOeoc8l9FuvErzkgGoqRJk5UdyeePkNLFmF2oUv8ZCW1XfCy2IbZSMur5h+RVAqyXRiPM0LT1
V3Ak/p2es3Krf6u2g2QK51hjpkas7uJ5lM6YcT2ZtuHvLT6o8Dio8UAL8qJBEtf3D8bW4qCmr04m
D6Xji3SNre8UNjjU7YKGc7O3FskEcDt59SzBGGAR3YCQwVE7k3bp1Zb2k7eK/TPj+LLWCaBFKl2U
sS664FRkMpzZZEO3TCnrZS4vWIHKHrjUAbV0+JeDIJKidgB9QK+19rYWo61U21m+oY0a/36n4YfY
cSB4B2/Bt0AIhHsi/vEvSj3DDf6va62MqBZ8LDxHgjjJejq+2Xrg4VZB1gIEtJQKDboYgU51/S2J
vbPntahOlKnp2/MWmsOEmHYONw4YEInMCjD62a57t9QHp+PbWdtWKaiQoUTAajsP3p0ZuRa/a6aL
AfcjNZHvHfWfKW/5yv4SbEv9rZI9mHnmmR8oGElZ9KNCcRaJ6wqtUuv7kR5MyI2c8Ia77qCeEK2t
eiYlNTlOrk6ltXqKvNJVojumGSxzFTV3y12yKj5Rr3OYwBrY8wQ/mg/2rnRDkSXvEigBt2pSXyRP
aQ532dVid2mnx7eb/Nm1erI7D/OTurS9SxTCtX84lk4WcasYAKgVM8m2R4BGH3QM4BGH2mW7art4
GNDeRBodIvNN1vpzEvsJa1XaVPq20TDEDgTSLE1N5NL+okjnnLbUcAJi3rlS6Y3+wrP6tg00zAJ4
QSRdzcpONzKTei/wIdI1dwPh2vvD2xs6Y4TIF1IlYlfUWEBeeBRGB9o3vLuYiGHE/R98SiI1/Kht
ZaIi4F+Dba14QUu/ccxNdUeHpaWbBGnM+iHUmesinnlnlDYqf/yyBFe0y7Pkc0hajFgjb+/qtJPa
LIIX9A455oPnlq+T3bBKL6kRStrllVvNbrHzAQltHvLJwnl4QtGop2+qnYQvTuxmtSSM20rzYRJ0
5z9TheY+N6UXWUqUIu7kGtshp37TWPtQUA3tWf0bXIFH1QQpouRlQtU0onWFNmotNajvRj8Xktvq
fE4IUycsUnZMCNOaBhGeB7CCbZPy3G3LSiD0X2VLzEjfZWXSPnD9gE7VZl28MDDAQ2eIFENPq2OQ
19qE7xxNMqVeHH8VzPusXzR38g4AcuTBBPPTCnc93g3SU3qScfcAtHZXIyiI6KtroOYs7JiBYTKI
qP0=
`pragma protect end_protected

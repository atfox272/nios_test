// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
R1nu+7Zw1uXvs4HyEccHPt1eC9BLEpKBR+Z0XalwmU4r8TsYsT6qt6za2MDtYrqJffpm6qYvbspX
k1b5NBiaX4FFmnEHuKzgONkb+vce1ODZb4vlH8A5RUeJ4EzUygiLnaaQ7fj9iDsnTkgKgWbshNJW
D9IKjQiKhBO/jLLMqPOnzSkECPp7YxiG0yt1Gmfid8X1esJTeW2dmgqft3usrRvxpWd/BBpel658
7awqqKHz0y1IIttr9NULbYtCgQnCbYNdlSdgqygD7oHioJnzITVbJGvHi2rUzkod5s6Z/lSkY0u3
pwb2k2nNjNck1IfKvsDyavwj7MyHUbNg+pb4Eg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14848)
UDvUQpHeS+MWviIxIxucqgRBdqF3VVU4IAuKDKFlYcVNhzWQYVw2vmHK7z8DBF8nD4ogU2iGn28R
z//gWMfTUTsTdT0gXzUwLU6kkSWI1dOFMN6Bn8G/ge4byzdLxsAccfspD1sVheO8c2urBXtGbxgn
zUBu6YykNbWDLejpPdNlgdYQ04V8X6OVEHf2L1VgixMC6kYaJ1E9arvnZhAF/dy8zaX0YihhgkCV
2q6J5bLswifW89Id2h8gPobIFewevb0uGSHM672Fenq6+FLFW9hKVif2Zidk+h4csp4R1xB5nTIE
G72YHq5Kwq6sEhXtY3MAMCvO3n5pCgSaERKwTl02hoW8dkVPgDyU9iY6wUr3JwhlbRsHWXB7KKmM
PGVgRQV5lVuIVuxNnv0sKeeHypBEgk24oSxOfxOl0pXhtHoj8D2KlqkdJ+i/L9LUELnxSwS6B2oc
XPysQv46xVOk5I5k5KbjeSB9pPoH6ZKToiy914J/q6w+N4Sl4hphrTV5SS0BdMXS/r81VuJRe56j
qmJamBJ8CCR2eO6m84BQAFUkx41fr9q0AnqMxsFpcTifYiqT+3E+z3dJ3iq5W2nM5AbgF8OxXfeY
L41gZLE+QEp7EXl5mDRp3+nMdHRu5+hKhoPmtxYeyH8zpxnPDKXUNQ/heePtEfRQzhotYOTcykhW
35bsp25N8+U2+9vH1JYIqYPtPf+XhCNGHtQPBJqhDiDmjSJssOYCPAfkNY4EXatTv3M334BH1+5t
5zGSumP/nEiJoWLnWS51dJ0nZ2PsQ1wVav4cMSaNRs9CUyN+4j2HUNZVRYBq5SxC1LegfZRTnp2i
ImpclhI3xUHeXfO6RU1ThFiz0tzatXvJU2rJibW3o+fpp5tpgULM3PdmMINvVX+5JEC0bH9Pr1gv
9p1E/Ijf+Pnep/folA1xH3ZYMptpw2XsnzVAPTnC5cR4NJeRhuzPuZQuIzHu6Hl+eCyTzATYQ6AR
PXTyEkwTskr89cO4lftljIvCZifRH20KLHJKo80I/hbGZkFgcBpwrRiA+bugdTGqMMS1DHH6U9O2
wkpRUf2cEI6MhGINxuW1T+MRluVvTv1fS2vvwVzhxOK0Cc12tROiAc+ACtZS4fsnX83wk72Qzi3l
XqUXyuwDhR7fP4xIRM/eEPzHGJCU3caHtuDjsqp/IUQTY1egtUsD9vKGMJ+sqcOfZb178aAdCLms
7yH5tOqSz9e8N32Hgia6ATYK6r9Ls1Zc3MPRijTojtNLjKdjX/I3IqLAt3/KCwnUVxF65udpe0ka
4qWrslaYweQbIBFyv+ofwJ/XZ/enbpmEYUY8KGLHPPepuAq8qy+j15foC/R0xjmUTQBzsHJV+2cp
1dbCma0duwTfep4/Pugv98cdSg+gltDwzolEsgQw4r8c0SlStMcJLEMbrRrlfxr4FMYL5Us3ee5c
SKbmzsGR1hkWL4rtQKfbBSiI3TFxusBO1gI/424PP5vgRvtchaEhnLyrbluEb9mWnItvmt9jvpTO
8MhDC/6Zd+Op64gIdeJAI+JXwBfgv0ZkSy74eNpAkBJqT7RMnjKVjzeQvaK4X1OopdXJ9GdIt9gK
QoXLviNY5rFH0rupkiHb299vdG+446uvNyluDzMP98Q9nmlKZD+f+jxZ0qSyUNccJ0ypweC5RivN
VGT4evxfqVgAS24yVfxAXXUeVG8eVG0hHvVXFkQEBWy/Aezg9oS2OXJjuoXWP3pUMaqDhIJvTIU/
P/SepbSp0rmfUdTn82fchN+/3ByyHXF0m1yQyvlJWNEyddsrbPgFcUr87EFW7qZXuImdx2pze61H
5Jd3uLoFay9f8Koj2t1/u6mWaZqJucRTu9uAhG7vI3Fc5f4je1ieWr+hVpiWYInzAlngzvzIZvbJ
xlf1bywJQC+O65JbVKvB4QbSaqscrucRna2tdCu6f4kKB8HfH0AnlCXsoXjcfw3vjYb1tNSn1JB1
q03OEMnVAwXmm6wfH6PxaXaB9nZl/OPXGfD8niJaWkIkCbc+V+/zc0KO4Z0oj6h/WO/Zd3meL31N
TcWNdooAYSGoV+BbZsP1LA9E+gaKhO+cO8hUXDGg+gXVfql1UyStDV9CU+HkDYwqqC6FSuH9y/Yf
gWeBB5GCXGd7Ud9dIwVtdqFKy935aqr+KtRdpHeJaOKhsMZqFYm+NlXCnsb8VYO0u54FIiWeidH0
2VPlNJUuDaqzpCBPHmUNZa1nEJkTBmpIOLSFGctkdovRhnurgkZ/rq7wEqsXT+5ZP4s7MFRvJgZo
cbK7PKDvKBY340eHWhr9T1q4v9NO9czqNWJcdXGj6C4ZNhjuHBt0ykaD/SMRTvRQunBfVPgedLx+
FJnWWsQXTK06hGm0QCSd/s+paYSvtynBELkJrhDdhrFDMb0jqZ0F5dhh55DXLYSLm2QkZhgxOZVE
EqEmpKI+Q+4Ha3CNBRFYOMO9M0A3ZjtNrdJx8RTrctEnqSlZDzJnX7MKHB6slOhHYwt/+6oYARnv
qQi7EalCsbnIBCpnpWHu8a2S4HnOcaptEVlxT8rUY1lyZF9a3ZzCLsSpVP5uM33XyQt7b0facBtM
RjarDy2hTWX8J62hO2r1qV9fr5cV/teJQAx6gNGwiTfUVltvsmL0IJtQPqzqLNoa5KVC5Ygl54Bi
eowjkJUSPYSeW4cfw0EkTjPUr6Ph+ap4zdfjPMuRtFK8F+QXTjuB5WeDu6eh0ujvWpBD/5q8X8sn
54pFs2sZcAwnkoV5ZHM3mv3jf6wLeHS6kvpeVF9jBBcO5Sp5nDONB9JiN5SQo/vq/hRBxaovRGzi
o3fcPAunYtDVySLh87t4vWHpcjtUovXV1u0X05SydrgRWXD6M35oYGudAMIVFLnLO0NznVyA+qpY
h1DLoWIFXVV2SL6/06TYHJ5uICnZON/Deq0pOejxofk+EDlmkCldd71CeoyTUzMenqjCkzJGSgZI
5OCrU3uRQh/YYg4p3/1nGsGnKzBOdg/jAemsH7rW2U3KfqGdTbD4Qk964ipMsnihtxhNLKVxozkU
7wLb7+mSVZpJEWDP3q2d2ruZYI1PLY4d5WvqqHsWDuQymjhEiiWnl+AyfRnrRKlwTAmXQdoHcGBp
mmepiifR++umEV055ZjsqbYhYzO4ZbYFFquEW+Vgpzc3FTVOOOLXHoOW0J/BG1Za1yYxG0hn6TQS
YqLklY3SqirNvvzCwxMbYFRFAgsSKjOjGeywGE2r2whm59ixZUf5HaDspYyzVLBNnJHE05zunk2B
q5JTIP0IQ53MbVx2ahTvKB+rRZLaip191R0emTSyMZeLFggkfO0+cAVyZ3xkHZNtHwvBTjUnGw0e
k6thSQRNhJ/uRyz6IRGGLiP5ZLgryaUZn0O6q36yXwWzrzkrXfUWybExDkNNZ2v5BCdq5wIgV79G
AAxhx1lY5NJ5dDd/x5LKqkQ48CgBpIAPT8Mb6991b3JqSpuxShnyjVYIer6v/Y7huRs6zRS9hAUe
2gPhk2JKHmZk8XL5HwHtCGf6oFNXaqHJOkwcl2wEZGJlrZj9EXn0rh58jYg9ICyrc7qds5RK9NZw
P50wof0j8EO4Qe/vMXD9O8wDeHYpnkIW+Fwt/S1OOGxy98ln/+1OdAqgAgi0E48y9f0Bmsp/ckFi
PpANEi/RlgY5NE+iMU1lYpkoQibv5weNhbEcpjDWmjUjZ+81WGEZPwOW9eqM9as0i32iw0T+DitK
kDiOhys2MSyrCXHeIiKAewb1CC66o54mrZPpY4+YIzMFOQVliACoWXZ/xV3djN650nVVTJgHhs9Y
kNVazD3Pn3ymsj3LmMvawnACMnpcS02Y8hP0ZrTGIlVO3bsfdtYk71R/nfRcxjfvaqQY3ofkn024
ajq2Bvvi0gciieH99UbfyufHe0fstZHo4SEMlmbDvegxq6wvhLqJeET5biVQbAdgTBRlHtzWO9Fn
IYLZ7GgHjI0xb6KW4RWmABcL6o+W613ZNSSN1f1Du2lLr8s7SJFUuDYI0n2Roef6JxyHjKjeY1RM
vpwYZ3HAezumEKkEV5uCFyYrSC4p8hhsDKOaYP3E9r+gBF96X9kEaxdhe/lpZC4pvU+PoM6IDmHe
7C5Ux919XzUygyH8vRaQPP0bqh8wZDwqV4ursGgXvh1eqtyogZDrMpJ5wzn54ZyK+8pjSz0QdhyK
FkpKyhiYie1jMQBNGafO9wuBVhSiQNVFLCqGbRFtKBk+8MmcP/p4haDFEVtNsXroOjYNcLL8ZviZ
UrYfACZriF27D2Jg4VJknScPI8K0qGRafzlprw7hvBn3MNP6BFyHD/MgE8WardLkUNZv2lRXn7Y6
VNlQPoRN3Q/yRqc4wGewpM7Tg4+6tY8v64aKhIaYemHDqRK7gQAtzUx8Xm1vseB16Xt0CyvyB1fR
2E/QxKw/0TN4iFFuzJgCRF82Z/V4fGe/6BihBPZ9IghSREfE+KJIC3vYQFAZ2G807GBAbepZsDsQ
YF4qryFrGfiKsvskqa8nduSk7pVHyCGFGS/dC0cAPUGyHDoPL0vvTbJkwafdEeuqRm2y4HeSP7JQ
rbGZBYA9C0v1kq5ozKmfpxq7dvZKQOtccnfHJTJspbYyy5IKi2qYesPxOKQOwd65zyGFdsUAs/Na
ztuuJkDwYDMY1XxZl/laPNYXE26D9ehTS7OZJf63JqLtklYCoKxz25QiGRva9mxty2NuqL3YgYpM
0GNN84iAUe5oB+RATs/KnibLH3qBRlshY+f12sFSZsUA4LX5L12pyK3hGV7lSVKHa1KvwTPouFPV
JCsVcjSBPxnTXKpGDQQoaKiwUZKGF392xKZDzrXcu+wzM/oaOxDLAQ1P9NUuM/djGPXRfsUeC8kc
dETN9BPqSG1SzkWuOwsEdFdqc03gKk8YAmFnLVpExgxLuHWtkogzDGrEU7Gbhk77fEWEkgAwi1DS
8hPIh6oDSaMrUz1G66V9VQp4t4Iot0NASJRUyNDoP2HX/3fdkcxT3/ki6ytmfWdEZSxp+MCF5NMj
ZaVk5MBSl6wUfLXtHXV+FXRTpviS/+yIxW+fWElXDadvfTjSV6Jlic5fK/841Y36PZ2USTL1C8I/
VgL9ofU2aDRHKOLJGnljmVwqaf4Vj8nOJEZ7ukSzPYsmQLFHrMzRWtYYlo6EkF3/zJGesmtx74Wh
iGj/uFI7neK4S7V7iwBE46KBIAK10ZNP6rLBlKS7585jaUJBUF0gq80covOFNc2F/jXCZpsmnrBM
kNWU7dEl23wUileBROhAl1j/S0ptPfjdWK7uaxV6d4FaunqymxxmD2OZdgSdkSg9xScjEJ6970Vo
fF3ko6PKSD7GM7OKanpsC17ELZZbiA8iPEvUrB0sBXXYwG/ib2p/quWdMxV9KG692shrq4Z1viyu
vLqbCErhLrsG6hOgFFYHSoBGshNyFIGH+QfQbmHKc+v24Hd5uUsJqulyjrNTY8h+SDBS5K5DIs3j
G4JxHcL8Z86IVrRcJujC9dkWWqDqfuSsRD+mK9DhuyK0zjNdoqBcolVvqeY7+y6SOC79hfQvl/kI
Ap3WoX8GHsNSlK3f0S4gnFZhJoEgvIVTKQM/qx58FzJk7uvlLow9YTEGHFcxftNJrOcH9N0yqgkF
lRoxlKMGchkDlFSMhppF9UAaM+O6aPcEJUKBoqIFgqV0gn8W70vEbJ9SkJuTrdZWELjii+4xC+kq
4q9V0f0yEJ1GSwc3uhXmIKMAN0ey3uTfc1XcPY4RWLY2sPGhIG4plp8dPrSUm5JIWomaeUh5wiAq
wpK2bZcjDwkDTbAlv6yquKQZsBZrfO2T+eCaF7j2ZzTVQZl58VUg5AB/cMoUmYmrYhSNrX7Ur0TN
wYq/Z+OKydHvxtTt3jmGgnP7D1rQR2Ha2bFDLQzuZi0LizDgCoP0L6U0mRm6BMMJ7x7uzAG4s7kS
g8tw0W1SBUe26u2EHLd9SfKvcXyRuNwh5qJmm2i2zdfyuC9iN1XNxM3gIj+tH2y7m7UKFIAfLVjm
ZZuQFY+pOvS+UCGiZXRFR5DNCikKGyr6RICAmHnAuLJosbqBLT3YNxPpntxWp1hHM6/d381mnJV/
QkwwdAoUlo0BNVChaYSeQmmJnI8U8UlioCvQZN5wdv1mtEk0Sz3gjDTjc6Lwk/ZwvJeyxdlkVVfg
gEdz2zWes+fDrPmOTasb/WB+4YzVZ21QLgQ82VRgF3P3BEQJea6N0eBaa5QPK4gbIMG0tjnDxAw4
uMildR5Rxya0tvhG2Fl9jAJQnA/8WtHE4lwapVhGxIrUSXtcbRkAxNxsTvTeYAoPf/EDbP9GaGau
U8MmP1jPE2qZylKWWL0UIY9g6xFpyIXwlynKExc9D3nBtuDz4EnjrcA2xW7mqeZ2MQPSONdwoYQQ
tcl6OVzIdlAaATXrWrzG4DHmSWqrqZmRLDxXVE24NeSNmXHQ0dl5T0jRS4wsK7tIGF/g9wamRBqH
Nfum/CDoEaFA1O9nLTEziToKV4AWTsmrl7SkP5C92clpc4YN9cm/hU8oh3pxLtiTrzDR1chCX4sp
26gksqK6tgDc83dRCQzcI2nQJUs7vCch7CjzIMzV3gKYieuzYyrlL7a7PCI4CLisFGrOHyJDQK1N
kW9c9NdKZcxAR5qoc5lmlynL2N1LTeb25iF+LFcCdD2cYthyhGTVXVj7g+ZHfOldHwVIYxY7abQX
JbqGE50lCxdUN1cXAA4ryfUaup99p7D2f0EtgCDMYHg/zf44TKE2YwTE0sLdTgusnaGmgDSoIr6d
TzvWSioMS6yHmuFw2+GbEY4jBc49gL5rHb7RAygaaH19rLxvR+8ldp5IvrC1fSoRDhfL8EGZea5H
nITIlL2zqfI2epWoFQ7LhvVUnJtz5Yfjm75ijV+5v6iyxKTxX7I2/SoDSpyM/H9Q4AWKsBamPMPS
qUNxshAL1plNuTuz08D/FUEBbHZG0jsIaf5v5IR31cbZ9KU7XyZmCA0/LVLbE3A2IlV0JV0cWI/Z
vxNlm7IurQkMo6hP+VoMVZuYA28JAYEHO/wUCdlBpZ9eiJzrRu36MTDOcHBjanwpOVpxh3A/KGgm
SbEvGXJpKWJtxyr6CCq6+yix3szcqp0SCKkNNhRKKTjDbV+EMPrA5qlr4uqs1BR2eoMwOOIs2+j1
FA5z1eUJ6l5TnaR7RSULcB6t+ZCGhO8pcdDcoU5GuLZ0CujSKMhBSxHwae3h98RqGWWSEW5evM8W
83bBS8AleELCzTcF/rTtLb8OZOpGGj09NiZBtnRBLaMPqaH/Al5yGY/MUH8j2m0jrQCbTKpswVVv
QSzvW0ou7F1kFTi7vlZByVQFU+gxjt7qYKFoUMfIZhmwdXhw7mCAPValY5K7wnVx0VuNwK1tsQ2T
TR2NdHI8bgOFJ2w7IDiV8JDCaKEVvTbDpcy1VJHg0K0LcIqSRCLq7EFzBMk6aM3vGdDcjF2+xfh4
fRpMM+UdhlmpuEivllLR1A0QoiVLvYh9rfT/oYzt6UE1M4q1TJzxbavNPE/i2WF/zbXVKrMhmNB5
4om9N11Q1qM3W+tqTxOjdOwlTmMlD/rGUYOd7oa4sJSIRDEosgNS8ahLhtwBxH2PXL28GwGG+A9t
e3no/xq890BD9/MWSiNy2xACIfC8mIwsTSw+oPYe/YowpXEQb70NH0Ls6k8d1GQdzvxRJEog4V/4
Id88P+gkP671kqwTen3qkJVYlhVMCZo87c0q/7VESHDKh/IOeEW0KjOQnVtN/FUsUkdG8tvAVGf8
YWUBZ18FcwKgXr6u5DkHHQR0s/AnrEcvhUpQt5w9HeMuwhg7q7X18TpPKuU5JOi1zbYMi2rKBYTu
tohYv7B0eIMMu8CbDjKkFI6lxmY/dU6olF9aGL+iCJzCzhYWrh0apuTGPisYoCOQSHN9aKpbg433
jjgCYaZnOWn1ERWudUXCYp6sV3HKPUEzRfmFP4oxt9WwhNN6GzVmEnIQxJImccZDfaEC7UfjV/eK
BxaY7ZnYwjYzmkSEkOdEAtudIV/hFpuTwos7r51uq4MuZXwHXPzfkSpZIH8Rxbllc7dzTC6PKVb6
sXQG+oU7+zrRZ6aBQFqnF+bISHyRL8VUxRZ6CCIy1/hOryoUaEFHXeqZeNAXRr579GqZG7cdJbdx
A394zI03RWEYo3VA6TmR7zf++ntr3l5gJaffqb52xfCJEHxk0y81qfT60ZhmGCnUj5ZehUex0oJH
mqWKjgKli+xhM/L0UoXP0pUZnd2uWXLnT5YmGkgLO1BPn8A+8VrNPsXp+ZcBrHWT6B6YZALOEYvz
xCtvFm7DgpVw3qilSxeSPcD8d7P9IBU/+W8X1rhzP+xSzAp8LzJcDWda9rISpeshS3bIHhxGqF7P
CjWCPjfHfaLfblzJrUWD79O6KtSGiDQvG2htmK7pK/g4OXgv9DUOMYpoZSIbfV4K3NtdqaLRniTD
nLsPqe0TCBjjsE5S886ezR+5Edlo8R76WpXpjz+doyn8bsjgmRnGci6xH9pA39Sk24cpqFFYmgyV
wr6uCrlsNPz4Cc1CuB4K2uHE2kggiOwKu72J+Q2LnJ9pwlyTWZjqpioCSoxWsNZY7lWSyj3RjJx5
kZF/RtA04mZQgsBvaEt3vR971XOuxBaszdQ999D+KeLmn9jHwexGztVUgMJLrfsebYTS3w6v/Gm7
oMvbR+tvq7A5yV/btXhdJ31WQeEoxZeLcdEXnqB+KMqra8xLQGB7bDFneX2VHfDq8TSOBoEdOd/I
FGrOhQEE7QXgDRwlnIP8VJjfWmVmiGWbyqP+XmJ0cHXunoThB2xn0XF59w85CvAvX3exJ33QI9Z6
9Yr8OBCRWEJdLF/K/JbtrH2vzffzdVqvAO97m3D+WPOtKkMOwNJOTkA+BfVHVO+H2gAHpg51o76Y
D/djMO5k9gPFb4SCy1cj8qaS9KcL80zghX71/T225OWHatBOV/M+fi3eoHxedej+at+gsC9dCZL9
fMnsM7nw83dIV4E5KhJirxOYDSBS6S7DMGeeF7la+pLGd8hHCW+jzFdbd2Uu6+1DXEGZmIjvALsR
VOyFWFYipAmrA5oRanT9VldksaRY14W3H8Ilj4r/FnZzeIAZ0hsG+L/dxuQZYmG8yt7mxS5bJH0A
TP0mTapJgHR2vffc53pJB/NsQ6tewtBpruLxby0PIB0Nj///aBAs3uSXNrW6QfW9XtxjUitupUZr
1sy7W4O5Jfgi1wkEkOs9OMEGFn68O4coXObS8hRJjzWJdWACx0nenGR3cUEAloslRbsMRzxAJ2EP
vsOR5S52jIE9iY0lDQ+h8+ZrZiSPa5UfmBocEcIim8QofCWxywRUfmZCsEYtune9auJtAjQIBV/B
jlzZ2j5gwxDOzyH3HOlZYTBqZI2rnM6z8XNyDeSKweJXLxqaYkmrlHVCeBR6O8GnYfjz4Rabs8Wf
as5B+ZrzVN27L6ozYQvV4mL4XBCS3xA+mTb2mCRPAu98eI7CGcwdcD2tSOz7HyRl9fqSf7hZD2yW
SR8Eo1Y7/yd8Flfp2iyrR09V7cMtg4/IPH8lhAYAuPyH9/OrflYgP5paOpdPsFODz4LigZfJCD2Z
2GsFUGtAO9xqE6Yy2pDGjK/zQG1WjieIX6rYA6/5LYKyJh/kzTF/FWxJvB1GbyQrClagJgt3fPyg
0KC8YC4F9g8MCDQmh/rT4vsNCpwKwXQ2Rux4lxTFEFwSgUD+caKcpfBQSjD6HvZFzRlXPaN+Op/D
7NUzkmxo07X/xshKeiZY0/B4SBfs6ZiqR5C/tmWMOjdvq69zFmsiEctn0DhR9/IrKwTEex4xHJwA
/0TWkSLmRlsRlRb3HtbTj8CHlNwzXiG2jjmoHSM4sNTXnuJuaFlRvtNJKqhVKZjF97erHss4IuBs
qQkp5T7TrIDoFlk/TxFu8Szr8fFIO6X9a1iFADi/UEXYhIkq9UVAVAJ/xzxbraTCUW232fHKWeFq
qLRc+u0aQoH08s92cMkEtZbd6PWmUIC6uv4yU1wi3nED5KkmYYqqc3WVpz0T4kTpAG7pAX056wqs
OCzDmEs8LrkHoD6Hd9cHxySuyJEGx0wVmEHNkIgQPfF+7LdAP4XwE0kcPFBGDqlLp4q/JmZqEzY7
ZT/ZPye0sAjS2HA0+wTUMSrUrzSAHM0zLoz3o8w3+I6E/zEJ4Y2GcT8ajQ1lOylkp03HmRixpkt+
2El+vNJd0wHmH1Jzh8pzlGoj5hAk2NWEjrXVSVy7rPIRswEgJmrq5x1j0e8Ab+O16Mm0l3jFL04l
rT8x2f2EiW017F8P4jwlb/+7XuCyhnfQeKwTehT88MZeyQWMGJhs7Z4i2IGe2mtKAW57vG/702Ly
HXgDedUnJwWyOJva6KJiaw52wdJKtTCFkyfjv8fApxaiyeOvFZ0ZcAObNBRMaz0MK1Z2LVzbSuwA
eY2xHHMWrrt6fpibjB69kOxachLgY2rPtZBSfqMsuaRNeCuGaU0YmWxaxMeH8FhnDP8oeCczbASz
8Zi7MunLXJwNm4NqFzbisadLBt0pCeaCvKVQt8xGbCVTEyWggwFxIdPpVm5Q2t49iIgeWcD+fWP9
lW53nO8qIHjYbu9oBUx6LGFtLgpHf+6kxVqbaQoXFhnkU4P2D7PAasejw+M77qitXN2j2DaOmX8U
uU1kSJwRZ3ou7SQZ9TDFZ7Sbz1y9nodkQpPMC2XjWZijmSlKzNpLbCY4hk9ohN4E10eCDhXkAarI
kSdzGT1o/gsukeckQ7gB3kERFzpttkSU3YAH1gWNngys82NDhAYCBrqcU1QKxnHWUadsq3wiKo8C
46VjKihO4yTidgWgzmhIE4ltCbaUqj8LdVwn27l7h7hin+rQskLvQcQtMuodBWr4SL3czet+komU
wnSduoGmxOxaVp2UgLnWUBnCTGJ/lK1byqvnDtYadZqlEpomlxO3NikGZtv4Cip3//5A9meHyoob
LLy8m7G7J5TrZiWQrewA+RpDsufN//Mfj4uq+ocCHE3EdfhvXCYJXUgNErpgqSXQNyEpY5zlSzKi
NJ6XKaYZi9PbYEui9E5t4aDmIqce3frm3M/sOeVNZuH0j5NrQmbxiWdKUXMioRSWvzYC529sbD46
w3pMxcNtiL04D93D5NASTZ8CXYN4S9S6BkBa6zOCJLlgBfPv01LLNRDToQ39lWfrLDwDP17NLmM8
b44/I5Kn0CleGSHDfh46xHe4lfmJPj5gTdnv+ZZR8X+9kJNlskZQmP3t2iEX69/f4abR5MnEOEYj
tz2qbenQuH4i6ibuWmM8zIIhn9/ie7Hfm6+2fY8ZJtQmfhldYcZ3EFA90u2iGqKg0yqunI7A/R17
dKrC/tmgX/GcCj6l09JqZSTShX0P668ozqi6HpaVYz/ZBGIgPIBH4fnsSuulCh6A4VcVRl0e7kih
fSxTFjYC7LtNmwDyby7bB1aXYZREZVtgxdai98n3/KABIgLZbWAhsSSvEfNiPRBxHRelLuXqEOtO
K0NRzY1IvjcatOxJbz3SP0kYx8WsgoTxrVpvpOIR6TBA5DlI44ZlUQicWhNSV+2NhpyiNY71Cw1t
wSdAfOeLX0hd1cv1EmMIAmNbUbw786Leb/OhS68h63eQ5qVoJp3MoxwXI5fY+vjnPtmVbyNnbE7p
N5j9sP43iIeb4L60k3kxHtENVYGA6b0IIJsE52aK87wLEGpKdZ4t9o80DRViy3DAvwWaeoD95a67
jLvWRIosaDkGjhneSoNkqUtFgA7sDCp/OiknhTs45L2GIbma1smUDwV7ayfKonyyUamBxmJkE3tv
Az4ewqECcRaTOwbe/rugeojSiafaD31eyKknw3N1U6R1NqlffuvhPLwsbTr76CR84kJfWu3PljpZ
p/5GmJqEo40qeAxSrx4e2bJc3LXfouEOaMwVprHC46vQ1f5HqCVB5JH/0SedK7Hu4oPr5V6tw1W5
y+fYXvrZwqiCwEVD1L/R0TfP/A3SSimRO97JqAehLHXmMGRkIuA2r7NRWXjG48UHttYuPj0RW0++
AyC1ojDpkUZKnis81HbwVLzOmA5V8tifmbRfdpR069/S+uGOSmZHKLPRuHyFki7Qi412VOok4mQ6
fJwTdnAkRaiMdrd054LneL5x2bqWTwq34E4RFXyHKhUA45fQPxaFzaig6GAsVFomGdMJusVqsvmL
JJ8Tscw8EjcaWx9gwI+SWINHWHxkXNRtitE4ia/W1nDhoWmRNQNWlWyv5OojuFyJkomQ/2XrjPz5
M1RzqnV8ETRYHmK5MBFOsckIYaz9zTzGluYlQvyfRps4BhsAa/tvKxgQXvVp5HnT+IWsCq82uo0p
mKrP/6KixljA1gSy7ykizHJfMNALTBk5BA2s9TBIE2dEU6nB+GHhiHhmZVipYbcQlXO863hcfM8Z
Ko79lWdUhJLgHkGLfJmDKfIfIqmPsz6AoQgf1SCdo9xvYZudZuIP3fBOHeKboQzzgQNfotitmG+P
tGIuk0sUA3BxQTkVgwFdsTMGCYklK2Xrh2Sv60x+mMytqg1c4HYWOctWD4Aq73L2sWQjD0PX/MyH
YiwWFvLCOyd2dTsA3VTRVrrHobDWG4kjpRQTI6rk82fEtE1dgXAGaSy7SJKepWPrq9WB3WhAjXhJ
52yWiKwgHWJ4QHiFtt9V8a+Vi7JGlgCb5s9GcGKiBz1I3lbRnB0NwE35DaZxaGyt7yQ0rxXNS0T5
svkBkZ/LMtmoLTJ2Lpq74+TK+Gl7PSvjLVowzNF5TjbJAT2oi0X9f76sdFnlm1cgmquRYCNFEMyu
iyjyBGwju7rhJ5b+ieQHGwhvjYfztXbb95DIYesxeWLN10KsNBnT+xYxD4PGG62WdiwAshHs+GSw
rA5nXaey3FJzzT+l1OT55YlmNT1nnndnLPsQ2yoPGxRC5tq2Rh4Rb3VUCL4JxLGlsJ47eeNpSvns
XDcUTADwqKYEW8PU1PoGuZhwgbadVOUPyDHYd+Nr6GlkypE8q8iOqLtXl3at1aaUNTMRDAtBV5RD
p7A06KUwHJA0WbUVf25Pd0TR5A94PAQVSFfHHNgtY6+0N6KhRmVIxtzL4++MACxjbT/3y/PRef+l
/qhgbgNt/g2zPx2d+YbA5y54hlgh9P1ilN5cHcAhz9AqPQuyWO44ADdCFQvtEexxhkqsDHlUwVZ6
cUAqHXfbkGNtXmb321TxC5niT76KPXfUVPulRq9GaKobN1BIZWaBNiLxcLUv/B8UwL46ZiHQLElY
m7KQX9NaZPvJ6sbhuidnccLIBLUklVlXx7GjH+xxGYmcSqVV0RFYfmYSWN/fRcV+VGvTTSUnUwqo
ZDrN92Dgn+ImtOpH+j/RSXM3911i5srXaCMRKGcJzBCwR/wT+fGu7/UCydKZ9a/TcCENbrIzAMie
U7YoQdil3T28JHIx2rM9kT6zizBuW2J2/XedtjoUWymfg5a38ubRkxpTcpgGyllqjhoP7XScmSZs
hG9Dp/N1L/WmH8R8J8t4yLrwNM3me58SwraFuduVY5/8nCS3oORcXnnwg4KOcCyRQzdeH+JICKb5
D5NUBfXSyT2G442Zb46rwx5G4GASANrxEaYUt24HbT2H5gDkv9frx1q+N5sQPKDq09JmDpPaw6nL
5/OaqHDt6141FMr6Of9xGjRiaISLsxjkhbn5SKZ8qAv6MFKvvDICr0HYFjCODaIkpbQ4zT9h2tVt
YwNn29LMvpiSvJpIov3Cf+1whD0GfmNdkXrV7yoe/Z4121pCsB0Dfc8zyIxt4hOVL/Q+mqlkPA/s
F3jTjF8v508tjWeyUG8swFXEgo/D6Q6Zde41pg0v9mRj2omxdH/n0LOzdc4HrApVVzqxRhRj9R+T
DOea3sFr7te6XaNe3qVguM0nkogNyYRTRp1WiHfCIbMDb5VnvW2e4RHwyq8g7R4SjL6lo8aqLJAz
Vojcw2ogbrtruf7cLx5tiXzn5HxiZrcX0A059AoVp/Vw4iSYnk45xVnh8PVb47IaTUlk9CBdnd9O
EBaFgGAQfw5lgZfbI8GPjk2ryT8WeBlb46yqX1xjElQn1G++D3fN/CJgSW4I0FiRyaUJJcDsGpzG
PrK/M3LoDze3AqP5OeQQZjcsTQHIYYOlX1P/TEx7pDXfTsHCFlTGm5iZ0zlvnyKZjFlzhIjwtc1v
D65I4Z0uG+kxEbyCPqlfx4RXqc7C2LESX7bTRuQxtg51lw1UgkvVsxjRy5FU4+l9WyFrl0YszoMf
zSDqwmSu1nghLENoPzhM0XbKT6Cb7SwlNq3JVI0W95fCKpFOuM6W3zRnsgPoSFFy2VvwZ1qxdzi+
rwzgT1QpWB7e0kSmj+vVYyAIQjPECfOokTLiaklKyy+dylI9YgfjjOoAdzW9nm03Nm20JxWqG/vc
Wbpok5LiWSU+cu6FvRQANi7emIBieWSWPC6oXuH+3VQsBlOq4GRKjHiN/dYsc+2SOiwwh/HlALHv
LZ2H2r8vMS15+ywsAa0mLLAT66lCqQ33tvM8RZJD7BzEm4trtood5JmR4gQ7FrysOHiw/AYmGi3j
eAF63LjJyL+5enxPqDxzi1ql35F8OGfgoHqV1Qum2seipcFwa2Hb/PwcXYwqFGlGVdf5Aohl4Os8
0AG3ixnJdXHlprucVY7DMB4cvhagdsberoZpNxUmexANr8Rcj3Rq66tUBPMBwoxrltkubhKIFj2D
yMBDHU35K79hIM8YPbL92Kd+8wopHLORVCl6B4ey+rspbAPpaLBNXgpCM5mn8UDt+qWQDC8t6d4G
Up1BVyZRv7Pt3POSnfVHkJ9dMUmBohwMnl0u5jVllQwxEhp9JciQ8dPNiMI7qxv9I+r05x8Pynql
Zzyr1hprupO5VERmpSOmJR17HDqNYec7U51S0lQhVRmrrDPVeZJ85sBsLao93yoxLUKwKVTjxdOI
orSMcjqGJckqSUxcT5gwTik+m4jsivc4T9Uw0T0LUh/hfEULOXzkkhnfPSsCcw/r+iLjd4gTZgvq
jp41Ve6f5+E+umSceT2Yign3xX5Gdg9cRIESE7VVLgVc81CFG/XeHgMBF5+Q/dnrbRqOUz2L/9Bc
4/jLqXDA6/0efrHAvaLFQiT4N04Rc8VanqzfrZgKhTzPugCkC+CzoVITJBtdng3d3B24YmqiONjF
osG/fxAu2n0nsCyMWdlIU/dGpEcMHJ7KH/WT83ZpvnO7QJBpS/xemAuakDXKHJ25uhYP/aBu01n3
iRUKuYw201q8VUSLR2EghxDG8m3UpOJH5lPYQHn3ISbubziJ9RJ9kDosJZuAgrML0BCHpprRb918
B1BotgTVY9X9kKXwAjy3UDLA9g4rZkzrGORpffqpkC/HTiuPhhfwb32Yhd4stobLWbxH/idzatEL
bg61js0Ek8MYEU7nCCYCQ2cPpEuYOZPe3vx9UlGla8EjlnaIX3dcRcBIP1tdTpJGXk1IPbGRZI2H
fOt/LMJOvIhQJ/ygOH+XquQ7Y9Q3DbA6GFV2q+iDrbQUIrxLgSZ5gZ07btN1dbGSkVK3uD25mV/G
Y4opDVk8ggMZpp3r0sgvXf5IKbEFiCkw/MOcLCK9NtiKowvtqyCLQF7QBSe/BO5EjLze6jf138Xj
3ztb6rcfXpAQQvh5/MD4NvjljRsUOGSNqFTfSwvqLw0DbNLHHWxCEwsT9W5bufyGgxG1mGJLyEtf
Fq82XpEhwsij0ou8szX5w+/sc/QdiN2lTqCsmpHmo+zJN7sra3udGYKGz+dKJC6mH0KPgaC1WVWJ
ZEXAuBVbxx9XNwcUmjho3lGEE9X8860bIK1qKGwrUCOII0LyZMvnOEYwHWNWTVH/xc+8Am3g4h8H
Stb24Djq8bNRQBka5iM3GM7aBooFwKkifuvTdnQQ6dcgA+YSpdbJuH75flrkWZL4osWWjxVXOPKL
3goHBgwK/kuAugVv6LF/5J/V+wJ2Gi4BOfUWRmHXslHEstRt85loLGdiBshAFDQkAJOb/zYPrLDM
5Ip7p6ilW4ev8spgI/nq1o9y2dHERmgQRskOv73lZ3vyXnPys8NgCWxEtaj2GOPRDQdcHLi2MzkY
xmE9w9gy4WH6oPcGPj3390k0IQ6aMSf1wqi06yVNNhmLhGrzLcMuBDHBATIu7jbA/cAdkJQ97mV3
S0/YKl4g8Jf4gM7QPUD9FGBE6QHjDPVbkLfQLB+RSn32Mm+R4gg1PHilbIrZTD/ghc8VhcyrW1RV
PFoo03iXYo1SXZoQiZWiu4n3j9BJaOORA4vKhOLjebrPDNVGToCqI4zLEnD81yU9H/RhALortnC6
blAQRB4KEFY930NQzgmVnYmtJBaCYtGfGWrjLFbyYiraHZVOrIonxAlL9cJsIzIMuA5psTQS6c01
RrZ0j6pf9zKkd/HY1QQ+SpCyrVt6Nd+BkVDTI4pRtvuigU1FfdsnFrJLckK0RgXOnjloSL5urefR
bGfkbk1GIDwyhOpgoRsh7WZ6dZnwsy6nvttuRBUmKWY2gz8lxvkM4Mrg75jVZze2o82RExA86CxV
3JSzK9jLUm64pnWTESj2F3yDBHB8vQCqYarM4AydzTAk8BCtTTOp+EOe7lrZsClyh9gYxMzT2VE7
RntITPoKncNCeQa8h3f2/tGTDwPJIJYMNXMcUsDivlucyHSv4a7CIj/1w3tS7mkiUyUZObQZiocf
gXf4FNWFInb+K2vTZzOx6oCHeRuqCXeZb5ArDDn2ny/B8LyxiXohW+uZb5BbaeLQ2B945AUKLTVy
zKbrDnOn5LFv8206Yp/UU1W805pViaQP32lcc34xwSIclYgjLnmqxOfqvkAVtsLIlyehS2hLX35X
HZlmGBGFbR286kfbiybaDJAlRMGjsWz2YA1Ab8y7thddyNpINCnR4tqgzbTfa08O0Mu/QZL/1gtk
Cyn3D6VnKkRfVyCL6A2qifrrYFuIvp2RkmmtD3s9qHQ573h69BuHZCt4jW8qbP7jWO6/E0vnBMKm
9kEH0BKZFoFPcpZI3rAqncZ7SAZUJXERXHjB3ilhi9CYefym4TjBX+fi9BD3Xi7MpbLJuxttLb/I
ipX8TbZyNVBs7OLUKmJ24FwJYnx+TuFERO+AUzMfBAFBs2zWB5tcA59fs+csEuYl4IE8Ui5Ucj2N
eAHO66qxPp08tP6/Nf1kH5TxRgx371QQhAF0I0h4NO/Tq1ksBh8T3DlpBGYgM5GWPtLZnPMIrjHO
QkJXTnQ3kQc2s/1E0M2uwHlNMBxNgZ54GhCCqmTzxcbpstTzse+yiTagfaiN9qUIOqbA9w0eei8U
6AmLi5Rtc+MmhLVAY0jD6k+IV3t1a7VBPRIEOkBWarXRRMFDxhW4gpAo88mVy0ir1QFzJYbWzUHz
IUcl+KjL02G0mH+2OIwbtDWqJnuLV80Gj2jJPJHi4ZXfuhzqNdygqt5QnfO1qfBogVPaRcdqWDOu
6DSUjf6wXtec9zdFPPlKDS7iHEQiyjiEls6nkCUJHYGZvBuC4U+FH4yl2M2FhEd3zR+ngNmpwrqT
O42x/5w+we0kztxfknYTuqdT/mI44klClHOBUHyuXKLpxWminMnvszY298bCdUmZa+yTeebvhuVA
BGRy123tWaywQ6doqEFgtxVoonx66hVauMidm9hoZkc5kAs96E18hbtw9Mw4W1oauPftBz4ss0xJ
sh5VfjgVkfD5ir7P7+jkdDcg1eyayB0iU8CNWLxhlkGIlMmMjEX5q1icFcPFII/HL9PY2JoFraxO
/pQCW1N9lkK8OAaPIScwG44iV6bDaHyZG+2MwDgSiOuYWamtMy/ioyQKH4ZHbAC37zXj7ERu1f8u
sZam4N6hDyIifWA0eBOB6ZxB+0wgaSAsCV3ygf8JmaWzsB5Af0CWdXjuFHApR7qYgswptDA5vBUR
LUInexHpxOM/LRjRMhXiP7W26Q+H0/02UPgAg6PuVV4+hZl1qFvKP+tFSgpy2Z5Oa782z4Keydbh
cFos4RpYaZS1NS5wJ+xcgeYdwQlsGjexBw4yjhXAs+OzsCJpKqWT++BI84IDjWkPPkOfDVBmTG3V
cyGSHrrAboLVLZXVPN0tl7GZ7SnH7Up3B1t4jhGWqCnSuD4yE0JVCsV/zAXVW+BCQyliCcfzth+8
hvbxzJoMmb71VrRAF8C1v7MiCCWjc9myIckH7tRFAQeUvznnIuMEiPA0RUXO81OvpVw6xob2aHRT
lrLucbR7OfpT8sHusRuO77iSm3EXfG3EDfaw94RM/RVdAh20NOG9PpRPFBfHTxqZktqwHHaju4bX
I3OKIH4b8mw0CkGz74p/3Zo3ZQFI27wCMNlLZbyVJYOZa2qoBYHdToZdNiGS521ym5RWcnowMKVG
wRzjWrut8oXYqsh12pJX5pBFAbI179+OhZYefvhn0G6pwBdGKWfse7rMdHsFee9A98+q//cNysrk
gO8/tgQVr2lxLdaDRLhc02wk38RkHlhasbhA6+YJrsQ6fwneGqWDtCOPn8Pn2hyt0QpcqIQxEUTi
jrQ/v3fBKOq3S7xgwkzoGCLNb7tGjOIkJmfjZt3xnEdjND8xfcqNqBFZgf2cwSOw/S3mWn8fVYFP
Tdi8EuZSUQxgeVgFyqim2brK+fy0hOIWY2HABx0xp7dkWgn5X7eV1IEBUqjIHDZdFEvNIDyFNTRD
JJX42R5+bRrbAQzVeP0nNrnvZsIlF0PWs3sOae/P3Sc+erkS24yrife8gY78RLcZO6aDe5jBu8+8
4x+vsobY+3pdCuciMo9Gu7pnXdfE1cyLy+ViBrSmBn+ig8UxEOx1SQH03DFXQa641S2XNOZpFnBW
YVY/R7oFKFYuX7XquP0wDFPo1O2gGPrblTUFwoGjZKFhIuVFSyky4FwBMX1O2L6bmTbl8bzR+9dP
dCAhjq25RBAFU2/2ejcHmR1LjopX2AvNrPGnSlgDKj7NcfQ1FKsnrgNCNXqPfKBgSHYzQqasN/Kb
tHnjv/906Zw/M5VLXJDVM6gnDdQbO0PVg4/Stf6UUjoMQJGycYzOnXW7LJIiiWo046qcs5JdJpSO
NPsZKrx1QXKyeIHDN1fBzcu1KoPHUtBMMXKhBGAc+UOB9fNLXjbq3Y90QrWLCALZWjtCyObNTQlT
3xkj5ozk72JPYhoC9n9uJO+I3/H59zUBI3lkR9Oly2vq0SMKG/SzbLEBHc06tM0fnIj5ZDScUlhQ
TABlacPoJThlkDtm5N2Iapv1o/tOoc5Fn8JhXTKKK6yP4M2+ZvgT8ujErVZ77yFyQZZSTo6ciD/M
k34LpTzSIVyEzBem1F1BxwgYbU3PG3F7zGxlFD1Os5+cPzuov9sAs3z23uAcbavpTX+D5vFnXq+h
DwopcQ5g3u5NlAlwoPpNkKgafDkN9N83VW8hXikPGaUlKRBqrNNgo6sSYRgG66f3kFrhR/dcg0lJ
d3Gk9dOOzbp5jzNvRl1iWTJdr0cZaMNyeZ6HVHs24HByONOzkZOZGl10vU136GFs/pmoJXIQqpAQ
PVeO12cFoch8Uj93CpfrWqhO4J+CwdUCCqqS8vh091hYcENlavTBrjB64xoLBEfZ3iGezwIlQbMZ
pDAiT0CpVfl8VkUtSLFnFjE8z12eoSxTEs4jAzWk6N9RNbbVGATmgXSLu2dWUa4F500ZSy1PzF09
qEtrMMFFvKmJbggQ8z0pVPNuq0pqiuz/pWHh6M78GfAvWYNwPSeKTtzScwviNrOAG8BIXtWKyCtE
4xx3D8QaQmkn8bmi2zQ/El7lxhRLf7Tqwmd8Rr9epDnMbYbNSWJJR2TFUV7i/9Lixjg2JscV9umV
5vHFLN1eKMaPjwHjmHDjoK9QnPSioIH7JCI+8g==
`pragma protect end_protected

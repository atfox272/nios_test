// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
EnWeBvpmE9n7EyK7oYu28gYUbVzIGR1hTqKpOysGk4aZVKqlN8eh5z+3EQX7CAb3gk/HIsD4ORUW
h6z7bnCoOMsoMiTNdjZ56gUF3htfCz1lr6PTKw9KaAuGWTPiL6tBX4R8Llr+kuIUpsskq2hbtBZV
1YnXQJlLu0UzVZ6+Fb3WMcriE6EqoGkwvM9w9QsfQRrkHJmSH+zlsr7Jp1hVwgwIYTmENz2yLaFk
zV3JoPhvdDpFIhq0cDzyrubStEYHpvM8UbD26kmKHhWC4nF2PFbBLYTFla7dO3h2cI4leSo1FmK3
fBig7IJabYzt1BNf4B7ovA50BCy5fJoa9s6Mnw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9136)
NKQeN+iSywxhAmxCGUlQ6Z+tHwIlXQ1m6TLO1JfgnzhdT3FQ9LqmWGc6tlNcgNrkP256cNNn077M
v1OuUxSjPtsa6J0NuYrkHC8NGnMAm8J4iiU6Rm7eJIEAmdA66WodktH5r9Y8kmXHO0bzQnoYux4+
LXT7FohXwDNdKneCV0/8pohLBoTQhTMFJ6ILurvHuuvmFupuVPNgVNnO9ftQsx7+cHcjtojoqXQQ
Ks6Ju9fgi7xbQ8NvuFAWdw0j4T8l7rWNY6Vy57siDIjTFw36VRhsocFnPKm45kFFeAXt3Aq2QpM9
uEmX2edXiUbNvy2rz4FPtsysQX3fD0sdLI5wRE9ZLg3IfEa8D4MUOjSyYzQ4L93iBJIZGxbpNRP3
zSZ+2tvPi85lrpAaTMuCsbjR++BK7J1K3/6B4H4SobTkPWTHyboaiKjkU8/daCMFqOQ/3LJF2Dv7
VM3bGNuaYaSUAdjgPEEJMwsmN/BukPVPnOKI75r5OaA4pwqSDTYG9JCek4HAYBLSC/Vd0VqbSIfv
d4LkYtpvwhOap3jtrYBuzXmNOcs5/VxdrPx+q9rKLh0DdRyoENPO7osPmgG/Vrz1+a6CgnWrqjWV
S//6jJHPK4t37/8ZdFI8hWNrgMozVyXYS15khKJffAC+mvt/6H45Z2w8E9u8wcL2UqONDORGrBHS
kRoEVUPadu/ESxkdDwnAPDtNe+FBKGMUczWHWXvEckwUE05inIyS2wIG6oIkxw48QUZUyNNZ5U9t
7lwdY+ALbUf9Vm8Pacu8K+LOOJO+xHOp86TD/IZKfaZj7CVaR2IM3Kfy5clDiBXKiXlELIbgJPzl
tvucwTcxmciCOpDFP0LJo+W+1vFXcaG7zWzlfrty4XdzS9DkDpQiJx6c/poVNOEeJhvqO5mHqNTT
C3gb0v1Ojyw3WJcsofGc/uU0IxbHbrZ80fl69Y4O2wV7esO6uazZkMfZsMekkc0lk3BmBPsFZ7L9
pbNKuD6vDk3q1tD/8C7+7QofdJR8y1lxfSp9q0KPJAFfNnJ0Nws71V0JD7oHIBSTd6eguaWEnm8O
2eEyUsKgkg71cOgaf9xIodhWZEmKV80SF1Sy+w3AkeNaIlICD0oO776U6Ua5qbhzobsJjf5pUp9Z
Fev3Ce+5S5fIasEAree6dJRZlizYIkjwObf+vwUG0M4RgZiwlc4bnLG9nJU5OoGy7pZmUUuVOzr7
bNN2SUZuYZ9HpZL/h/KylTSzmpAdPj6qKqgzkzVNL6tDu1cRLvl0y1dJNoCgJI/bhGzDZGbwroTP
edYHV/VSw0f9LZhPh/ajbs02LBXDKPI+hgPjPAM8pfXJd8DKpFCKokOCzm8eFlsj9UELR4LrIken
ZXHcq71TiBQVb4oiVKwWw+He98bdUX5OsKKxftHMKpXJds6CpfrVmb1scKlgX+HQzyDVpYBQCEd6
gjFu6ALqX8Kh1ZeYKO+uNEXFpbuBrIL1k0cpOh6U+07fqgg+0U+r6JSHu+wnWNwVI3Vc/v67mdYE
9LMfG9Kg1KmUBxRhdwWb+JFFRG+2ngQXde6Bavl8uYF8K8Fv97maI0MGOb66mj1Dy2b2h2Neop+M
mwJF77/JyuvWX07K2hm6ss4K8smH6a2IE7EyUC+xILV8GP55MbXP69Bg373TZypIiYguvM2wT+c9
kvcaZmHRkdXSk1mAaWAo17JuSQL9BFzhnrQf4T4g6hyzrAwOgfxmMm5+GEJJlZauRkOhZ39RVRLx
W4TsuYgwxCeAjc3QZZxx9M2qc7CaSpEQLtaa+yrO5xepc5BxkwkSNOlHYeDfs2xin/n5/ebXN+iu
LyvYqwfpHPZbCsIdFGDkA5tLV3fTlP/ypoJ3OJXlctMzgfTIbaWCeiP8YKNOSLema6WTBGrRzbMQ
R6Bxu1Uf/iUK0ZAEMQYZS4IAlvWi0rLtv8ghNdli01j+7warU66AzxxNfQE21VQEKOYTBX8Yb0Md
QrH8x521p/a94nUZoJLNDafKZLpDilew9SdbzPUnvWugx45Xbyo26Y5ZRMIVdc+mXGG36HZOORAZ
efUSjzegoE3xnCd7iqPdA69HfSJ1/PS6lLhT0rp1Q+RHr8FgKHj1CAC2wlzf5Zz+KehCdVBv0TMI
ext2qll/FZkvxJ/hyfZSl/9fYPLPG3wsg48/7NVrnTarnl1pmQ7k2Jc06hBQ71pjug6y5gnRqE7U
ByBm33oZtmnYB6mawb7wYhuCkXh1ETOzUzIFTaXDHFpMJV+NuGxGeZj4f5nxakDuPXPNbLeLi82u
I/szKc/FF3vT4laGQlDViNsiIiUFLvRoZkjcSdpQvz3A3GIIX3FgswjmqLwSXPwtBIVtSpK3hd4e
JZm9TcVseKyLWoroWnqDkGhDqVkqH+aB6gP3dLhGctyKAdZ2Ol656xa+fP8cylRQl9l0IpJJRdBs
ypo1HbgZHAADmrmNdeO618ab6QTh6+j8rUB2QNCOuZGfsRKDIOgYYDtprZ7VkudGLEaNH89d9tYr
xwi/w5iBtSudLGWDo1YBYbhA0+Jggx/QDCyyNpEblEjv9FO+Uhp0AgXU/oekswEz86CW9vHwxo4R
Dwc1ne9WeK519PWY4c00tdCvR9FCYOJWdNjjvSA5mq9YAp9kw1e+ZyO+V3uxnXp5oUIyMqvMICP4
WQ2U/GThU6BYmWWZbVm9KII8H7tN5yY7jNO8gduWXlsHFAxWTZV6PCd8Bz4Z719A4BsrKmPtGmsx
bHQPZ6AJOXtonNnSUnVWzW9zV+aFfngBbz6p5i3NIw7QQVbn9ND17klHCaFvtYp8Q+X3l6B7Mst2
KmYI3/elH6Fsk9iajT30gWO50+yJJYMf7xkH0FxWbb1OnU7k3zyNOdl5AYztovhZGSYpmfAIACWg
6xApnprCLZZdN+ahM1KjVAeNVHJBt0vlJGr5Y0dbVh/FTC25362yJRTb6mEbqoRq1ajvw3Vlwkga
s/YWEEmasuTFC1CY04CgT3/6fK/79a6D4n0BlJKBim1lrSHf67oXfDi8l/C1xH9YIS4duDlP+y5I
ud+6B/ZiaG8MR2h+cxHe6BpQmDcMPfh+KRkv+aIk7af1asXN29Lv6FaA15DRJNLEH70iQMN5nPSf
qXhSse1Y4oZSJX06qtp4X7ypVkSlIxMRtUcG6fabo6DX0EFz2GjiBybqDZfF1CnwW97fFJop/BVq
rOBD/FSQtp4/GGlchtGaU5jzXTQp6zSOfi1YL6Z3Irh2TGXAofTbzVjAOgJOOekQjFPggOlmGtqL
xkqClSU5PnMLybI1/SiAMAzL2/YA7k8JUVhokAzzDLyLZuoiEVsZKPpRlGsVYg8CcBEiBHOt9JBa
XFO+jI9kSOowKmaIsxOLWQmPgJ+13NkCV3XZgwGV+LcIQWMKrArFgPaTTRwHLTiC6OnJo2Gy0i1V
kyZt/XLGM69d6zOM6nkjYYLH5ogyRnaKFTcOhu+IiYv2kpRIa3LKWLzv+SCXs8Rfq799UEmFMqyQ
iartesT9C5Exwt4uwBcSE/4hQ6AsdYqSt3IDatyBPSw0AV6jAADt+gjVIQHq2Rzi27iDMSL8DW7P
2PFRQ1X6EmzNcQkfVtltyn+knktjfYpYUeu+dwCILlNfoRwXJkb8OQ/hkfTbHPQUrx5gFmSeGiY/
1BMlt2RnzbBeTG8pfv8CAffh3eOz2VdFn3vi9wFKL89sk0UGJSoBsPkCAAHZJgntt4gCJbH5+B88
2+C+kqFOF7xpb4bJxdUww0srF06/qrx8VtfZW7v5yd8dbMH8+MTTLFqPPT5VLs9ndrFrYwI+BcXE
2WI1+Iz3IixUqdGk9hgCHMZaUETFqP7zMNID67JlOlNfvaw7jp6vw/2AIHEdRJtys9R24RlM/vcv
hEOdqTX0hrX7d3epF6oyjTS29GeLd7SJ2imdo05RAT14spf0zglLF+W+lOkJPN2Casi+CNeLumwf
UeR+2sKs3Nj/ahC+Q3sDsbPtQLiBSJ5ynhmN0iikvzQPO1Fxw1fbqTWzNxazWGG2tVCkAtI7rNkE
kYhBJJvbMITq4BKuIwQgFciwpqSK5gZa32OUGEgOoHNZqHvbLc1PS3Ha9dil8yYdMR8xLl9ayPy6
2rtGJNTNAumP01ses9a0bmUozk/svICEiTGjjZpTGjsaehMzeMY3D+BOw6955moX/Kbi7tIcB5mN
YRizv1NJnABb4N10Rgm36fT+kCV7JpFLGBZObWEybebnfWcjtBfpBi2iCD2E8vmvE09T4QEgC0wX
5vmv8S5onHSJzQgx/RTkWMU03RCB2pxGVcMPABTD2DsouDmlRPNPFCuhGRWn8rb36O5xNrITR/vv
ou6Zv9H/Ksr2DK6dr1AoY1EqI5pSdMjlCFG+HAAqAP6UkyLpo0DnjdBPO6PlJctzoxILR9Hou5Xw
gs2zHrupHTMZ0FMzddNJDKRoWmEBE+Jz0QotRUP1YRDuGWvmvHEhjkmp0vFAArkpDmxCbyUqNQPy
rStHkoJ2kHvA0Lt9kn6cRtt3wc+tylq6KczBw8K8xDxo9KhKKBLabZq9H69T5ERW+Eps8j6YXjPi
PYHlGpJx2+XvUwoQ9c1GwHkYO7Gpks5HtSEN6/1JKNcU/Fi0fZOoqhnCPnZVGKuqkrm8YMnKXImZ
50bkAayqLEAfTfdyKT9xt2Qk3H5jl1EoKTfanPU3EzRTNQqSy1H3Lh2aCOoBPaYpmPV9AADQSoUb
fWSwmYIxqJxpbxmmCBM1oxbYotrnbqGcoodqovLBY2Fj1Rtwq3E66NyDDkar9ksTUk/XIL9rxIty
J52ydvFSILaQNDbLh25o1qZFkVOzbPB4WxKNutfKTf8AArxzCK6lBOMaBZul02X4r1KSl3t+t0bV
wK9L2Cp0A28Hi5olLhuC5iqcsZ/yE/+kdRqkaMvzkRyC05RNM9ULXvprwUEVui9RrNRmkExIpkrc
TdVFMMOFvk1E1lHKh9LbN/GBU6uzzzNxYw1dda/7zMqANehXoNLN4pieFe+8qC5SXNqXbez+rqbL
tK1KhWjjy8btnQZXQ41Z5LM9L2ZqarRmuQK8gEaZgSfxCJyMxUyEYpeJoks/ubxP0lKCOO64TNCm
gJo27WDlonK/iNUWLP7BbRyDthbK42eoh8seugc5+YMptaeKsSe/AiWb3D/kudfV/p1PjZVBwS9F
XqM8tTBanvXSvoOUBiruLv8OgY1lFGzWPdfaeCDLZRK0f5pkUk8zf7rIcUawdDdx7OFwzVBv4NrM
NKr1joCT4J6HqeHD+VJeIjLU8xAGRIj+Pr91XuFnS9hQFrWk+yiv8Q6MyFazOJyCC1H4pplLqv5Z
VAS5ilaWPbF1azLMVBLkoaYHtJ7f2RhKZdSd2W8QEMrHCRTVK1/n+imLCANWNHtA9pXzBqRVSR0v
tGoQzwKTpNoNHKjy6Hx4I7nIBJddSnwEfJ5fMtKFrtg3bvJZzS/4Mqfe6fkmUtUzd9PIASU9G8IF
ERfnGwbTWnl1oalgOxkuylM+E6gHo2aE8n66p8tIcuTfNY4ITc8/LnUFtCxLkxUvqE2rK+v+deHC
7QgmVgX3Ji59MZqjP+EhnAU59UGx7/qFcRQlGYjA47ginBbGPw3q2NO5wGfQ9R/iYfv5DAk0XBjm
+DLbhbkethUajBQBIG2PaMo65z3jmI6utAU3FHKxSd/pI4Rusqb2/Wt4Wnd2gmukaQSXc3SW0O/t
HpwtmVlv75UHYfvs6jf3vZFkL4ZK5Mv4LIuYvy9IMWw0+sLbdK2QHjOkDu7K/ZeEpTpGjshHXK2o
lrvUTgqnJvzIdJDKndro8ylj7aSPO54A5C8PjhUTQ2N6GRTHL1mVRbZQnA1Z9yVi008QfS/n1Q3/
AG0ErUXRlIgYvw1yENL3zeTsxL5gpW3vO7CZjNOnEHtGt8LlxfyROKX05gDx9alEFtiB+6rLP2ai
CBo+u7Wj/Goim3m4ic3/h33Zu7Iel1u4bxuq3/BU0YIeYiV8WbBl0GvUfawKvYqTy2I3S+PKP2J6
VpHwP+xzxWnP8MOICiR+mb2vGQSOnoJkzZ209CR1XpBgpHOgw5dkLvHvedCA6VzYifTNEpFGf+ND
SF9+2qNnqqcv7cHlTuaZVYIPLG/5yvAS2kw8cCsrE8L9w8vgfJi89kj6DJrAy9+BvoUcqiO2fuyG
mbPD2ferh/n3/lJ2qRbPcDvHocM9L5NKCeXhRPIzH5BNdyPKOfn6iVm++1RUJ2NsrG2DUUThg9qi
C5xfnOJOZV574frc9McJi4diiykdbGd3N7XWKHwHloIXOvcRyC/MUP2+Ju8Jbtix9Y7cqYaNMglR
kekYhI9tLVAGvc6EEnynnFyzI3oCwd9/2gSn3Fbg9QTmG2eVwoQVBlxoqcyr6L6oV7n9KtIvtGS1
nloX/HmxPDzg3+nqHMXRGqwMWnWna/9yiILzqb9syyD13za2Hnn1Im3Jx+f5rhBpUtWS0Wi0QArZ
DCtYi/BewFpo9EvxQewg7CZWXIyVvh5v4FQbRaDfTQ7XFWqqy1JBbBnDfQaHlIdewRhi7u9krUWd
lPcHli1VMfSiEAGkUUpKvv+0APmYX7JTf0M7BK4Gk1vERgd8Mfuutm0fU+HiOxnM/znab0X5Pvbc
7h1YMFdG7tcAGF+Nc9ySWyCVcOWWXTp5KZsDqN/Tk6DQEHr4gbwWBbqVdpxGw71QIam6vmaltirU
0vFQ83WrQ1i9BOmuhuUAij84pvZv68cXc9gjZOAaBCQAGO/ozSQFUXAXnFrNl2XeoyezgA+8jF7X
GCBgQQB0sOvFNetUWIq80i1bvMgcmU4O5AJg7GiwpiZcO04TQUwgCjWidDkkdxzvIXMHUSb9f8am
CTKNNJz7dj21hoeybmyj0oSXWtkU+QxQgYU+Kq7amgMW5RBxDnpzUBEU0xkA9d/azxWsO0nmfKW3
YpYVRfFbuWRyMJ00qjZcwy2wFh828q9IbgULJimxb5gVCaMRXHkDrkkfAWVRxoxP+YQt56xZFmHF
1ulzxEwMBP6wOmJeGLwaiUNiZLTSxW/Q19jFOg3c0Nl4RceCMDb97A4SdULeQSTInINeDG4kwhp+
XThVMIII5rd5X2pfQfq8VhiwW/mP2q4mMjAa6uEE6K9Mr2PQSl90g6E0z/plRrl4Pr1nAnQrgBfw
fsPsYibzudsfqGlgXIBZuDn7WTvIM3KjEY3i1CNwE1a9F/kpPEUOvBF/VpHNXXpyY1GQJ7nImgq4
p/1nUD9RWjFjp4NOKtZ2T5EQ1xoBWPDZAdUTzB6wB6YfXEW6RuTA3fbp4eXs8PsOJzfJ8Qu2xWXJ
CBAnHfq2OCUcS8B4xfwhv2JjbW2mx6JyeGtpSRoZluSdzY6/ORcV7fX1HOgP0D60coMwPPni9sib
WKTF1swQLLAANT9+QTS3HvDQ1FzruxypdJhFGoC4X7UaqjSoVWNkpzX2YJbZKGoOwL2sz+rhlWi0
V2Nu8lb9/VYqT+x2MZ7/vmtJU84KPgE7WILOj+ThFSthkOMdA6QlqjuSmI+23rtfRJjKScaIr9My
oI+V2xDJPXy/gYyeLwekeFDj6PLODsug4kJNVyk4L1XNkTXCmBpGCbrZL3jq3/UHgy2wa57I1mgM
Vex600XGzxtSCla6XMg8RfF+S9LcRytRlRAiabF8i4otcL4K+5dcvvhwfSEICxOcR0FeukD9lw91
jfP8GYULJkhhGgXsbkPeUvoA4TTw4YYxrBU7c+3XW/bpCHqyFh2vGy09Mw3P0PaSE5X6uUGUd4Mw
Kd8rbSEe1r4IHCOr9Eyow7j1E9QtLLHUMzTC4n8PBdu4/OmEs8Vy8EjPY89Su14zCwDRTkTOxptO
DUTwI8DkSXhGrKOiuP8eLsTbXCoNoufXnDhOLDp4XEhV4mxckNLI11cYIuCA1K1Py6SQPp2sqMDv
N5TViuFF4bE5rIXhH0jkHgfefX0gES4YjBVHo5B0p+2baLLjSEsE3FMgaB2cOw01VRnhmzgFP7Dr
Hc1WtRSyVrsROo+sSboxpTJVIpqkT6k4XvNXT7BmPgqtyHV8tAHKkDKVFV3fOZdzdRTf3CoJj02O
XV3zp7Zd4CvFh0Ndpy71tZRcseTitLvI9toYKxvavgTYPGt3yeNW7hr2y9loQpq8gp5QbM29ohrR
81GleSfTJuySCiRdSNbpGLn87koYwnaGrSkKbxCIHO8K6Iv88B3WeCCD/Z8EouLrxJ9xVjWh+/Nl
hTAGGWCOA2OnlM5wDPF0456B1Qa9q9brkceN+S9vcq9T6j/5sU8J5QGVmOtp7BIUlzk2F51eO3vw
IPdeX2vICkuRKth2M52OoJ81jZgaBetGv0CyzQecsguObVA3SN+uqwTrp881id1mOXPFWFAlUdrg
Qgg6qqaTI/XJ7T1TrL7zQ859Oem9koAAzT7IfMRITt6K/nE92R19kbHOkzbCgSWQt1AN22ooWodg
oXTG+X2Fh6EDQ4M5et6gwAqD18XjUL0elfgN8JTTVROe1qKNKnZyZ/pAL3JgKRjY7G5V9FK8WH7j
GsX3ELWPfTeuNL9avE4fuiu/EQCy/cOHzhglIBtGJMt6pAfUCjbEHneLomlYMsL9j2jHkTS7hBAQ
XwWAM7/SDGWy6V8/9MluTf+gzI6tqOG8fMIODiCO3Wj5cb3I0n32qkC9NT2yRX3S7gkHdCvpgSgD
XL2CFokOfsvGqbvPBp4fC7OSa8udSlz8/Rp6IDTEKiOEjyOzs8UmqGLbyKCVO8Ty8BRa8aQZzksH
cKyel9N37mEpdwtVAzNisGRpGMkN8QkNHYDwhKejCbeLCyb0rpnu2ldMw8VkrOL4/oytFszQ7tIg
JrPPJx3MXCgc0FDjJUWBAtcwfDlRldPc5onCDB476VCAXKzqwjW8MNK8i6TbmgTnC13w5QKIIqKg
J+0QALgyh+Pvqbi3+JIC6GWqat3Y5zW0oDZDkmWAkT3p3EPaUQnrbh5nfu0g2NCJn0QR2VqdtX7l
NqlnrlrgiKIcC7w+c2iXI85HrjIf2wmJpEMawrJ4cbsJ/P3saIKjGWOUClTFI0AetOJtuLbR/qzw
4iwtvIIwaNFg9riQhOc5aErd+1EJuwKqoTN0KIyyoEwd9/gggdte9eATXDBUCf2508CtxHTxzkKc
F+veqK24kbclsxtrFv3WChwynbWrnIuZE8EMQDLg/aYDS+tOTHzQ1e0/rB52/9nGuvXmX72tzEe0
VEWmZ5DM0BTzZEMQh5jvLCgXNpZpordaNIA6/aF0ooWVFMtGxzf+MjmP24vPC4ZaDeKvESqAGUoG
f30BE1+grcQ256LnvRisHMKSoq428QQ8dD83TcZpqom0f6dCeGc1GYh0jhzRUFJmGJhqBAt1rsKh
SchN07JXAIUN7oBs4sFi+E3BI1MdoAm1s3q1gINGDhxAJAwzQaPpovDDKK8ekYMgDD0XkoDy6bGB
1v2dBk9NyHlgFsXw23kWr0mHAlLC0FgMUGy6spPVCtdky9EO/Hz7T8W+RechSzuzu2xeVgHdykyl
PSsXefcBVCQWNLdOJhgWYCRQ9y58Ddu+op1gcxMWBuSi8S2JguuvjEfmHfTonuqdBvf7DBCwgNKs
C5lZEabmZVilVbT+iEUvxxKdwqE54eQNLhDzeNlt+11PmT+4yeldXJ2sZFVtrzR9VhGG7n2dlzhF
7Phj/cbO+XeXkV++bjwUtqUi1RIql00gSceG+P7h37QhytVmf7QaKhJkuHz2YDYcuSWjyuomAqht
JQAZKWj81Ekq4t2BmMfe7IqiDmqUudA2Y40qk0VMadjQN2cx/lmtWpHDM+fW29vPkl9TSxq3ezz9
otg9EvvWktLx4D7yfbzN5DHCckLA0yyiqRnLBLKFIVxqXgoCzKSNE9RdISimXA3Q0NKmRU2tQJio
IHtA+6uFP2/setfAHzcwIBYRXv2JZpX53aAZm8Jt6637MApQ16bDk2BUnJMZI1zgp0qrGob6/hHz
biZ5D70ANTynPZ7ILSWtCgqcZ8kHLnJBK9LlbCX/YdHEWUDem9r5ve13sIacVI46ywAqup453B97
NsLn2FwsJBdx0Qhxs8m94WSsB+porn2fCEHy5bPk5j86bQjsjtc9Qc2mmh0nspuTTuuEe16zaTw2
p8UDwvSK33Ua1cbLwC6dqhECGG1Xnb3b44k0SoEt3MzsCoD89Q71V74+dYstQIqTIy5SNhcurv9A
SsRfUSUI9M3UDZQPrqp/RKbqoMdeDnVGTBgm32oh06CUNQxGI9jFP1+Jl/NFJeHKlnvBvYbq1g8E
iFl9W7zMOdX8cqEbEAkE4zKE5bWQHPx9Jr8f8BirEPsat5QjJjV7HbEoYu0wt47bqXqMytXfN5FS
4FcafJLZX4VSBcFAbsAhRnbIGnJdpfaqDZvftxOXWXlQ9r6TwMBrXze2CAoyVRWgmWkObq4j/sKk
Hw4sHNBy7oQlw5sItie1wFoIEY9l+7X/nqEhpnnpOTSLbPhTRfWpWdKknko85Uf5omyMDu2yx3t1
jKS1AokVr1FxqoSeZLFJJJTP1HuqIJTAubjnqw8BO6j20KRfA/HmcxZMnPfJrlmpdJyPvNUUPa6k
4NuqwmfrscSODfljpsvbJwzNy58lV3GhTY83xn0x2nzzm3EMAfFTOvmLEkWMh2Q33nqe3kurJ2oj
1xGgeKeRjg4pqth9SJGt6bCBLL3/R+JPLLIR2hv766Jo1bXA9VtiC2cjbf9mZxiHnBoAqTClqDDi
zGURagzY5cuQM3lWCgQik2Efe5/hywgnqRlyiVoBhrh8TXGhj4XeXGXPkmPirO/imBT+qyNh6yzx
0IR33UbS+F8Ip2Nrx4ez2JSo9fkWpdeY2XbhUexvaq9ytSOFHCfe7K1ouLFLI2ES4S8X/bZ+C114
JaMBJHb87JBlscEU6n2epN86v6E5KZkAH2Qti1ZOx96lPFiexAhvhx5e9rpMHYB751i/QqIsCW0/
cRxYqT/otmlQ3C3BTfpiuIygh1snfLeuAocWu3PUqsAYYi/lFTLcq93hpGdVeTW1ZCzoUVEeysvX
1JzV18LsuObu2bsgMCfX1z+yk/KHPB4Dci6yZcu8aDACXYQam6n3uXRXdBbNUiyNZ2r4oVzG+zPS
VvcSV1sNbr+DreivaIFaBvP+unNppdvU7dW8rio9boKObs64isLJL/aAZgoKpv66YQsUU8K8/Yg+
NY4nU1ztfVhv/WuCtqSeDi5sG97PHggFEOUe+YV8UuFz3PGLpbQh4ZHNYaonHcdO+XMJccFY0cHG
S9sBXBjkBxQeqHIiZKPoaZrpMHmUbv21Li6fHLvqKQ8z3Eu89SPi8OWf7ChK/NKOVwgjxnc4DK25
DkVJrryPmCgeK2EcRxA8Vc1RyU9J3R0D0AyLtTUJqdhHhrbXLSSGwIPchGrK+fbAP8XxLGN73GcJ
mNEZQx0vKM+HY899/GGcdQJyE1oFWKZ+dwdqOMfixXVK70L8axSz8bLZjv0CDKlivZZws7nq7PR+
2dTWtrfoPaIFa9NrGeWDfOyTwRYinSP02MutXC5qRGahSrtWhob9us5/YwC0AAMokM/P5WuNA0zE
aQU0sHXriveDQuBm65q+qCLVN4daTTHOXHMq16YhqCl2wcydRsuuCG6Ds3wHf+GH79TuF5pFsJan
DrRbhL2fqP1xCF1kDeGbiUdyl+CBDfhDhR2agBv2fl1p0RsQD7qTS9GPqcUNyduOBbE0NEYcqG9r
o8Ztvz1vW54S+yy2C4+N4n9zx/Su1JdoiXYOJns6a/TLUPcQSUNlsSRA3gr3aOhCcQemRAagKujD
vxD2/ekDNxKzRwi5gxOWu9Dhmd7N4kAZ4/BuKIlkbRk2ut6dHuGwKIv05i4/eEDdhTYUUMITC9OA
q7jG2Ub+rz2bWDbX65MoifON7eco44WUN282KdKmMMAY9MjtdLFzrXXBk1VPUgA59NiU60rvmFJZ
+RHt/yT8mLIXU9z+U6j2SXz1yxFotvgYiHXpJXQldZDChDYZGMD+dF+KHmRnekdhgFC4D2zpBG13
Zn690Nrml1X1qwHMKk51ESe1J0DwcOzDF5kUU4QkfKVu4T1Z9ybVGWGwZ4uIycX2RkJBm6HhCTwX
CrK+q6EG4ENZM7pXke/kTAZ4QdyPxaM0EBtzYmmfTy3cxK8V+9KOM8nD6KuUww/S7S13KrRJ7hgm
Za/QDMQ/qu5zx9qbiaHh2g==
`pragma protect end_protected

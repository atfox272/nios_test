// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
yfxVBk5gSywd7i1aANwB151HmgibC81ghAFAP7BQD6Y8qJNvyX3i3eNW8dPXlq6Arhx00Z9s/Owj
mPAkjWcK/TdHiPSzfMvpdxd5OCa2evbnnQLbQ2IS5Ts4Gxa5Mp7dfQDsLg84TCaJZcwNBPiq11K5
G29vLlXECeG3K0FokcSALoYPzQLpVstg4YJwpJUFEIPBchB/5pNHiPQWdAC/G3q3DnTOT0WNY86E
nTBP1vRrjXiyMu8vjtAPoIPib+2TkeM1dRo/cPO99yukNZBCsoshReGFlYcZAEkQU/uu+71H2XnY
LI3NLI+dKdt50gTUzYAtSqOLx0Plr00EoPCXAg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6256)
2OwLmVvNpIuTKn7FWB2Wc7EMs07UKxxteBDEYRvR3KIxjD6eKN8bmqfYZG2cpeQ55xcmpv2zpI7v
MJGUmKKpOjZIywnvYSyTqU0u91AW7kV8KT3NsQ1LRw2nRaYCp0Ek3wwpQM7SUXzexm6fASUb194O
I/yqLnpZOEzsMAnjAa10af/cnicwpaX58wYJguGc+H9QVwlbGm6cQo/Qx7cL1AOp2cnDZDhLbKvW
cl5+mcip8lEQjMy0SxwPDPV+vUl++xBOvb8V6sWe8cGgid+MhgfNdOIWpo8jtWXQFMCmxQxC+ln0
QGIS0eRdkVnzSHbc+JEmVg5MIFDhJwkHNkha3mzrShsFNLeyYhciniIVSn8DepJAdrSfUPhKbWN9
m+fmU1bOqGgCqYAnI+7Hqv2SAEJrEL+C9YV2rAvUkQCwrF6R/OBHpLcSOcsFZE3+RQrrLxy80TX2
uqA2sOa9UIjg8xwp+d7xLpZf4EQXIBCpURM6TqZFIJCojvfFVymqvIs6sJDOFANddCtix1r1a/z9
zdhlx05iidr9aO3vqwYXy6qyReyQEDrzlis14jq2i1zjlpHpLtT5PvbBE/mt2jwWg1w76avOgf1G
FRULJcy2Xa4cDaFtp9CcEg/w/bB96X2RS2btkIri0+GVEkvgukAULomiM7crJwU8QwrvL2AOlyXb
fCX5EB7NX26K7QpjgcqRxDws0bnrrME8iniCCc3GH0spX6Pp+PL4IbAoq/cGpkQA6pg4JBQcWz6y
7A2TckzhD6XeIIDsaOSiGKuTZA2QMJDJWYz0t4dsW1ki8dYmcl2jRtJ0bZTWorpKSyrQac1XYAuX
+5sBHFK7Cl8cZCnlgsaiSKBHnBHZsnXvjkam9sFmuSbiRflunxUheFnvF4Z1uDKKAjd4pM0o+Wva
ghg+/lWOjhvVc5Ohbz/aBFBn2i2fHJzmL3lyAt5BPnEfamkidI0KMYw4ZTnKBXZwRCPULZvOwCjE
zu/XErIH49fbB4f2lNYlrkzFWtW24ysEC52/vsguAT0unMDn+wrtbkixZyZxClKHgXHxHngM+QFa
e/y9OFf0kkOYmuAYATsIdmr0sKPf69owA1WTYU3hMnMX3zHcJmme6JDGotwSXp7fjGVuHVmIH5dg
nI2xTKulQf1KXVPMTxGsksMWOLFzGNKMHbTdMjywerIFFDumMjgfMjLvixeXNtPGhgs9YBvScf5D
P6PZIjejVytBdm0MjgKDinkKDH8K1IuaHcy5tJH2MmqMdGrB08Fj++YCRdkQfJ61a+3eOJtwyxHn
Bb/CG+u8yX7CdNnuNRm4yo/QbTfLuPjY4IDVDHzs4qiJy/K6c8dbuFj6ANjzlcA5f1WtwcaUtjQZ
iE29cTbWOwFS9NPgAAYRhoE69ZzZ7wpa/fRPkHlBPztYonfxkwP9eotgNfNw8vQNgFlps8P7mzLV
emAjOZ4av+VOh8Wv6YLnCOhCYM/08FR4v22jXZXeoqlxBVVjDqk8ff1cZQflRA7B5LLiKXABI0ja
1s2tI3ThedkEKgJJWMipkzH9FJhZ8szSzO1eQQPnNZHS6+zNKNR/+Ql5OQJTDlqL3MGGDB82UHKi
dF7KusMyU/Rj/kMiEg3nDsmv/DTVXybdjs5EGYneYM3hc+2H4hz9coF7j6Tt8MHr1FlhtJC8jHhT
L1NaRYjq9NblVXmLsIvVFHh167PNAvw+Eqej69TR1ij5pEjin7Df0f9IH3BIe8B5uL0am6vkqUP8
9mWfwkC8DxPVLKMI95RlNbE58v7W1DjHiX/s1MTDmuDn3fM71FBX2pUorhcsq8GuFV8hXTYcE9bp
zyximv2BrqeM8UReSzdQmC5lkqRvsd13QhC+HSkj19hUanxJ9Hc6j1oECiH/yv2mElQyvavtHYdJ
cVtJI0nVYvfni+zCyt7fg7CSQCBepMxglEXHgoPo0TtOxy4inbOJHKKsBflWtOWPCdM9P0UIy4Ct
WzgE9M1VWo9HrBLxgAuOb85CB05nqJRc41EcAanFsxJ6sLQq8q1oSJcvc/UM+nodVkfCKxKY6ZoZ
Mnv6Yh2xJQSjp0ImZc3DWUA/WyDHN4NhjzqwpyWEkGR/+LQd2enLNeWgcjhjK0QqayCOAcbBDjqW
9XqjoCSzSmyzhLfxb0nlsm52H6A3Sk8Irrl9raOupebfma5uz7/LzK0MXnFH8N9jFy9M5t5F7jIq
cMgvR0e2V/py8NzITD8ABM+69bHzgF/NanflzWOQz+8lAS+M3pqs3aODEEM9skucyMUUX14vFLSD
Yc0wv+e9pIJmDlQjxCVW409eER8LeoVgFX1C/ZYsme/6Pjkop89tDF7VOqcRNEsQXtR9NQLSsi+h
s8OArAULKfb0tXhrGHfWUFRzs4HyqOrt4EMWbHEh7c4SAjRfirflCBeFnIV5/pdPz1QoDQgxXZB0
P5u0HHe27drbCGhnlUXWFOH2F2q3Z5wGQWgKot4e8mPmAcvht9NFhcC/ILUauUMgnI5rXcfQRfmZ
JX+37NbzYd1o5SXk1QK+BFRIAhNB+HOb2B4wobrQYZ2dZNxHWsUFT9PgEyi1JpOcLXAmyEtBiVFN
gZcvGWOu7t0JAVXaLtuEyNN3SQlslZSHPOO9sUCM8wVo1x+r654XjLALoRhCPMltWOuQKbiP54i/
VrlYqc6xfL3cztxldEeejCyv+8cZy++U6mAN01yeHTBEFCsbu1SlZfXUgEfsBzXwGIlPR0zvBQtZ
ghJ0ekmFeuxzrR1RwFJwcqjSNvARYcdApnqFLgV7Do1ojVzbSur5EWNgy2YQTcgSq0QNeOmHkZzE
Qsvmjse9k2vdKlnnbDNv8LgLg8tr/YecbMgxkL49fs5zE7Fp3QKtMunGKniZuVhuHZvsIj8Kvecr
krUFxIrIIIodN8/yzOqift0D1FgQd4+YF1lnTjLl4iJNjAVK47+BvIektxWq5I38CaBUWSyNVqnL
Z4h+mqswrTi+I+QCLTI1m9/ZPJdG71jIQU7Se2POTbKPy5Icsp9k6Rzlx6u2IFgFdqv78GuT+2EM
12MQU/NlkXA9w1KM3R7m7ehdie9mmkVkmcSjiU1hcghMVOp/Uydn65EM4IgMBZ1NAn+adv8AH2XD
SJuyCvEd9ZjDhIgBUDNke9u8zgITg4z7ZzBf5hrRAGBJUs53uqc0qqFhXoEv1pqAGsg6m7n1Pl43
r1P2+vIuV9U/4OI5hd2KoQAyD9PDGr8pyfblA2Zlti9s7LB+FS2Ob/UaQ7aBbOSaq3BdQiyFI9cz
1TDhGlCTv2whf3Hhfy5/sOJ3Rr1DvLZ3qHmWk6XLjG+RwE8YvSk7skxPmVBzgwHnRLoI1pIrXPfL
IihMRTL4PIRpA+K2X9at6W+Di1q36TVs0j2uhjHHura2ni/qFG/S7yMkMq9qGS8t9fASrqcGxOWh
RlW8OIzx/SrJfOQUXauTqdfgM+diVhwaRkKMe0c7ikoshk28QnUtnb0daDu917Xx5+xMNm75WkOa
05vusJjlNSnGpHZhdcArA7axqY/KSuyQGCgZZTx27izSSvG9JCxgcT2Eqi0olW4vrjVZUX1PvXre
KML8+y+JducC3Ax3I9TZ5dG7XbP5uLEl57G9/tSvbIv2GwQc1cdvN/1xz2tSXKRhrRWR9st7zBAk
ffMNO1oapaV+yUL33/oJX2IqaO4pClwGt9wt/I9WHNdtQF5XKY7IlVP+Mm7WNOZGP0EOnaedsoYW
Tf9vPOA1mQQN2eFnkY3PRhzGGphuF6M5xOaIwWrUoNqDgVuF2bBOISUZ4ppYgfLOO+byz6/f5MEV
9Im6XnDufej4A9kErzFjI362athLZIhm/XJHZWfEGLQ9hwWosv3uZarHL66ALrYS5yF7NjBVWnPw
KITQF5kQJP0VJMCozuJHjoTznC98Qtr4sQu5lfokuKJEx9+WywWfccT+Uo2TaX4mhrXclWZVVVSG
/WvK/y7nemlANEmItqsoihbVm8/iDqfzi4S+Ov6gtYDG6N9YgrMrGriGThfhx6tzV/HRr0+a9N0r
hBZZGCpUWwkV5DwGMg1olbwXRBSuu1JR+DPMjgblQ2JSbscNgayjfsTvspkWS1WTeZhopk6UzhhE
b/quHI2LW6ca+/7QtKWxSubrZwz3I84BTlhwGDG8kfgDc0oBLHzqZXJCYd5EPyTEbbOYBWkUqT/1
3pREmx7jzTKRC4sb158xjAYYUrJPB8DvZ6ac5X75M3aMPkQ1b1tAeMe4ASwckyKEA0Y3FiLThAVt
lMYnrHMBgoRB++qyn4FSfonCkSx3TaezWTDZPgur9PGR0LmsmseCJNfLautTcvv2fhwdVFGuyYRh
SJct2bsXCNaWyALsOkGF3dgQ6zdPO0l9d1Pa5GIedIxRrO5WGaIFHyBCseyBUbULdOZZAWxQxVQT
G26P8e9NFb0FOnxynRAp21Idam6AjXEf/oZN5hZND93sT5w4x2tZvnW5z+vywCQ1a5L9DSJlKd51
NEhn4j/NbMLJYoqU5qCwPRLV0b8gVPE4EafsSWyjuySuBh4w+KuuloG1SMWVa9kOOyJdGpUCPIQT
6zMKOqeBLSWlgj615OargkqsAENLqHNBeTPcs1YW2KQX5TDdUIWvdbWEVt9v7s+5CAGdlEu6J0vM
81rhaX1enRCBaY3W7eQH46xZilf0gOh6UhFNntwsP9xM0H9nxrYtzDLz8vx4HaLTnvO/WMgeL/bB
vNVbetnd8Uif7UE2o6DyfdJO0tCLw1v8gI35858AnVqvJOvVbzXro2Qz6daeqtySJQ2ZuViSJ+H0
poAisgDSaTNsqoZgG8KYs6Jt2pcdyTo59HG8MCT3CvH7h8SkhIhfnuTl7MP3BX6kfDu/hlUzyoL9
VSc6wKd6M6QVdSC6/SRAuwO8UxgkKTJvoGy92rIWsWLQINomjYczz3MXiE7+OxJz+sOSE+QuI0In
q3T9BBxtsZu5gIaIzidkGXOG7TwOa5Ew4koUeFF9AeP3Pu4/k6gtwknG/5ylyQ3DvFutknpwuTnj
CqcrNQl6h0nQtEfZ8OKpbUOwZqa1PZoebccwsfDCPnciLxkcdeyldZvMTSpdB6vke1LdyHVWOZzS
aNQxzNNUgY4EjZEOAhjZbjj3EvJHozCnZ007mKLohw7CqnRLghwGrPobbtur3yGVLD6Gdivw9zz4
pbZu/VFmaWgkZ2oKeTYU0tdo9q+Shx3AM6upFpl3plOYaUahHZYq/khS1fpJnp5OSflnz2MH56kh
qh6asFceSKRYY5+2yGvhwygg6ChMvVNZBS8vdH/VWtrvVJtRL2lMhYbaX5bJAIItwU3ivwCbMhoR
CIACggBz2Qq+Px1bO7XMa0T3ticTZQoprogpkb1opfRJ+jAIkHv415qPOrPZkHjTRCOM7e5fTv8y
FXid6ckmmttTnL46+OQZ/JfnS2Sf1vLUBNlJxZNgB7wDyg9q7+B3W7vCZiJHk8+b9U71kXQ6R26z
btwnSqkord4Ahv+BWr53RvlXjniEkuNGP04I8U0PoJShf2eF9DnmgXW2Lq66GpSYA+kPdHtdzI6Z
MK0DLL56NQ1G/dWjT8nePokMy7uwfGSXmshkogpnwZ10ROSrwBPXR9mYZY9MuUZDtQGkGkwglktQ
G1i1v1e4UBFLNvQ4FbgGdlsteojS8+q4J7bzM1my6TnvN+t1JyoJ6q7BOfFDHzZp2usJRBInipzN
7WQRY1cyU5ZhGY45d7P2KvH26TO8CWQDGAoiVTb4AL++hM6pQ2P5pLgJzvOwkMeZqetT3fVs7Eyl
q+9uk4I8Cl/5V/UFlMm0XQ5AdjSBBSKAcW/lesRgb6H1PTwSHnN94VNXZEW4PvJvYtlbvq+bfbrE
Hxzqdi/dxka9geiIfSYSNloPjySdsHUMdAEIRRHEM0HNMnv5PC4UYBC8yES/2iFbjwXhD5SD3DQs
QLdGAWzfBGl2DT+ZGp8ytl1ijZ6ZXLn0rTM/YPF/UxwB+hf4yw4Pk0wIklQM3zVpVcrxgA8/ZZxK
UD5Y0lR/820GlTMSlJV6oLVtKj11dEq2dKs5xoHotGbzQZIhp7eRo9Ai129uj+cc5iAS4EHfUrvm
k8U1u9YMHH0be07a67TXiqGYrWZJVNUpeWTnJbYqNe2g3a/FC8DlEUf6+HxoMN/JcWM5XaMMvou4
ydcTKnKI/mrC6c0RN2qr5ABhOwJ11WBvHzDPpbyu5Y/cyiMh+szczi30M6zIyeQ01h/1fGopKETn
b6W93BTyIatklFwwBybNJKIH2YgoC9bqpHAfQoqh2Pzzp2G785S7kiUQhvSKwT88ZJwirkO2JeyI
IXLMutHfyh82eFrXWGKENNcZrWcJX8fGC2VRwBDFXRPY+Qr7AcLh4yzj8hTVmvNhBo3x3l2D7hw/
WDzsTouwyRXFmt1sGJK0ama6BXD2NK6uaZtMkEvzi5RvrwXR9gFtQ9spVP5j3mSH38rPtED+zILk
wLRKiJcydmfz6PmJb4t86M5MkdU83For/9imPCHsyxATMysaNczLB1lJuy/ysyoZVvEJzRdVFi4U
QMtnurnHkJakGKZeVLs0zM9+uSf+p9DcvJ1cnG2X3gN5RQtT6GY0mvAuj4nw9/CcZJ5gWENFXgru
BuUU9wgZnyBfNXdRDppJeOyO1lj4OcK8pF8ZLSFlgn8tebJu63l1TjStedM/WJbEqJ64DRxxlJ9z
ZbCyywyDmqi/gMofN4wVYTv1TCgSiy1OAWB2QGmv0SRIqVEawm0rjG1hCMvwPbgHINKE2Y8myTnj
Sqn8VOjTbXZqdLgG7ezL79k3SsuJkFaX8XDTvJzUYcBdOFrxTkXcBWseztM6IeF7uombrg1puHjw
Aaqo2KjKYJ+SpZjJlVBkZP3nVova7fh58MnSmKHi/9GFDgfcL3gmEvs1esQjIgM2mZ2e30HUAK59
LvegfEwri/6rqRgpzIbtWxRa0Q5OVumT39Z1wQSzX7KG/Wk/DmwmdYUkjkroHCdORJcQwmy8m7v9
s85VvHdcngvoSSQYMY2KDQfaskYUAXC4vjMNA1PW0Hree27S4jcncc4fh0DCdoneuB75zfK0bSuI
lkBjF3dws+vmCCeDJHbLwGjXPETivfl3pML7mZp8U6EFxnyw/Qf+O8RYjDcSR3+IMt5ZcNfhFPba
pyLW5+Ph5eq20AqbiOX5R+lagATLdgKxhMxlerRwn0Aq3S/+WJLbvKpSzMA1l6mVbyyOuH15GcuV
8U3pQLAo8C97BBXrIX0wdKgYMf61Csg4L6qFs3cjopOyl0YyPHb60S6kBn8ryxHDbH70KTOe114l
+tB7H/YO0GZLH4QD+eeZngvYpvH4fztfqWIvBaS/urluW1g3bozO2Z/P6Abo2EpgbhMnBc9SZT+I
Uta0BSnHZOpS2ksAFU5kyjJBgNUWpPqaoUxvwOgLi+vHhdTfZGP03gngcVDXpHoS5dBE3tyt/DLQ
aRElCIJckIMD7mr4Tq390X4un6NN57Z0Bvs8yoxDMULAvuGU5nTIojyEQTSLBZTpwm9rewxb6YOn
6ZsIoSirkMjWCOTbZm0QACCFJlgVVDRNl4lTMvK6IVK1SJvC3Yp+AkN90FQT2M1Byhg5Xy4+/qVK
EionPq0UaQtAsxeTPZ2JmupKlfeodcM1IKmyx2Plv54YvS4GWMn8v2lQtYhnoM5MWkxO4KaijbCT
Xe/i7A2LKeHyAe8/JGSAFvTW15SMFU5JGeWUiVcYDOgCmYUdiit+Zt4PtYRrVpO1I6cuMyjxhXhG
FZLXk+3wVDEnltS9dYojtbTiCwvzP9QDwHNqOaExdTOXEHbAAoLKUP3iUYYDzaOdnM1fYuMBsg8I
DH77K0TyTMpNd50dcr2re0kuiUfPNbu/IKLZrGj7ggiqrzUKG4m98K4cf3OHr66xylVqj/5hNoOd
dV5qDNkT2tDzezwL3LhBXfK1LRwekuZwhb9eqckqGA+m71FZIRFO2TOLKdRCz/VMCmt778l4d1OV
ZtNLKdeNYJKJhJbhkznla8voYzLmaxvCpQyYiHSosm6Qi73nok060uo4IQuKcaJcHfJsafqgMFyK
QTB9WnLmbMMAH3WikWyxXI3+CGOqsy0jvE2mNsSGy15r/h9NiToNBp0GIUT0ygHdFeoz+dM9dSci
shEJMI1Pv8I+7W6wC4FKPoeBSrTXxHEwYNcV8H4kVKD9rmgyXxo4mRMQNLnUfbiV+ifaXNF56ZsG
MiQETJmI6gBUSgwGIwNBgKfHLjHkKwU7FmHG6JevzK3d3Glyf7xf6Qp3CYieP5nKnzFQmVXaNWyV
tIKULv51hVvi9YBy2bOcYnkv59wmnSkDxMZwm1cLuDUNFGSxlnpSPBL87A==
`pragma protect end_protected

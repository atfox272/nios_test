// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
M76viMRq2ugugq/5Tyc8xQLN3YHtU7+Cze6AQdooZV7oC3aTpbpnhVS7ege3f4DTfvMY0ZDMj34p
jgsl88leQ08KutKhtcnjzyYMlxLbLseujnr3YK5srLCY5BTfgAqIeYeZh2LZtTeF4nTxGtadVuB1
MiiNlQrZFzNhXcy8T1cqU47YbFPZ8IXI2MCWj55b0qvOC2QDNDlXtOhARAaJuSF1dJdhjwfvX2NP
8LjVkBqOzvzcp/7LqSW5g44Q8/xHblsG10+OoSesUYp+QxC/MC5rp+nh5S5zsGoq13FqIfi4ueG7
7LojSl9dln1FcLnzE6wX2QC6HpTRgdz5MoFwzQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 24000)
DH1AtKi69wemaWjO1/rLEtr6ciAA4LRUZKU8s43OwVSapoIXD1So+R7DZ17/7l/el3bGBSkl2EzF
ygB2Nw0gAaIOol/iHh0wE5gmYdG2WutlYdtcD71ep8/ZF6q8nqMMDRLoOZ7GGVipK2moHv8ktqgh
O13sgCBx3V0vrx2Dc9BOYCR9iDhFpHDFrdikiGFIbWH1yF9nkD+qeovu2BTqoNvDoByUWeB9G3Uk
OvgB6Lw8qqyVYJpmbGQ098FNhWuo9+puhpnEnCKgC+82EpEFK63IQy/CusESJF8g0Z5bnB6MxDWV
0itxwuWyIz6eehssXy5Fg5G3NgQsv7VSZfW6vkrO59mn9NFkPyOfBTQhL8DkjGR1u2SXcCNyZBOB
FypwxDbAgfVNWYia6awoy4Hv4PwMNSvwGKPoHU8Ve5ekfZkBo/wNxc28u59y/e/drdwU4db9blv9
VM0MuKVj9KZfQR9sLZ6/ingXYLWulK7cvKha8wQHsn7Bb9ShVq78xGFAMqacQdfZ6jReeTiCQ3EL
5a++P2wF5iXqnzWfVNZp9mEV/kV4l0nx4hneBUz8b/mmxKOhffjTJeGj2dX0lKYf8jr7sSA3YoQ+
xYMPko/+gffLhTc7+IODBzk7jWBk+M9aPWuzXgV52DC+9lyIlQU7IKxa1mPtEqElW/kpVnXMmCHQ
aUesk5wsQxmTzS0Kr7vRuBenwMFChvVPOLk03VJp0iqjYkSSveK5KJqyXvKDR/Mjo6xJiG7fDbjP
xmB7FsEe+6Gg5YaTVElGhc0yKZYfCYwFfTnaRXRQt02SXcK7F3FQlmqVpIT6dU+a6eISnZi7LyUn
LgKg59Yebb6Nn/5iNNgzUnHC94TFase582OubVTnpdqdFsMePWmMx15X90wRWDYPV6H96c666dTF
ZA4lhjdyC0BRW7sgl+kplKtjDjQ1J1XqXAE87k5yZjumofFraNCLPYhDWNykfftDEejZ8TxyTYf0
BS9lDydIXYx5ugIEt+5kTPCWikr8TqwIycoF85+2aMKpD2ZGCs5ak/to6/pWT7cDrpI2rdEiqWuI
NrkgemGQasdJIIy4R0JufnB3POrzylyGYD4Wzw8At/v76o3pRrsTr6qobq90RPKDCjeUNHwwUCAG
YTLcCezeSsmFC+0d/mIQieHBZWc5T/G+oEQsuJmAAIuND7JzeUlxuz7ETKz8nrZdbpKnGu8OQXSl
sf2Qrp0KngnJ5YlLCFMAJoAoQgy4v7Q2X2EbPxKlc7ZHaG/6u7ZLrbN8SAkhkQ1ZhFP7Mc6GSzQ6
XHzLuH5bkzz5OqiFwDjrr6xvAyOw13umLIiM3aBoApJzTasjLtghPcNpEfjjF/ylySqhyKqihAOU
DwT4L/lhp/3kkO1JB1sgwKcLfoJEtZ4ocEbGIR+zimxcCDtx8MWc+A48tisOu3fK7vjpSZwj8xsP
GDob7GKawbunvf4Ybnh9NAiJCnFhPWAev3lfrW1K/8vf2aGn0BKIrRIkP4WLXfZax82/Y/j5hZ5k
S1C9CenLOXZazGHgDwjQ7PQ7M3xb3X0HlG/2uWAjkKJYgsKiU6uZ0YMTyABxw+z6MD/ph6tOcN70
y78k3i4CC2uRQKSjGUuJ3S4aDTxrxQgADhuS5KfGbrzFaDpa48OM6Hs3CZPh+Q88JWT9uFL0FOep
bDDQhN06y6Jwr9XP6WXXV3MPfd8K2MpE1Ti597Yb79Ce7o/64OQYPMlfJ0N9rDoX/R+QfVVPU/44
K6pGJzkHmSg+ylLQRAw9qUXIS0BMOdWVHDG9RPf2Utsfs9E4OpFn+UC4lizmM+/XiqpcF1skVjwm
W+HrAXw8jMiXHlHwCtTXDSdrwBsvS7vmgsLGM/L4T1A3MUGeohWepsw2AOn2RJ/TL8o2OpKMKWtu
nh3P7jTgfbphdBHS20v1iQQ/7O0OHpwazmC53jmjTCj3WfvYu+9YhXOUw9KRZb02qEhnW2EP6VnE
8cv4utVPM1rEl0eBu1ctasN/phQ0wK5lVSL1Fx9sEeq8deapRY9CFysulrr3M4c4tyAnOQeAlAnM
sTC7TieZ/CjPbR0KG2V7tkIzN0CjjkIdFeBnFAlWuqyCOjSTnrKqVLHFwheIrjFYAzeY/y0B/f9B
E4raSyTrUeaap/KIP0OhxjsVYtHJSmmkUYbJtEWmL0Ug9rxPniGvL2iJihScl7Xd4c7xZAISJCOV
G1PyYtIqKtIE4IUa0/C+y2us0lHkB3HqqZtnM+wggX4JVyq3sangOCMbMxcmkbenfV/UsQ659r1X
qek5nvd/OiRoYt1LmvbUQjBatTWBW02AgpARGc9KydtTAJlzCq1QPT0gkiCxsymEgAKJWJiJEXnB
73Ffrkvq36Zj27bQIoJAw3FWnkFQADl2G3PMQUonyO8wTpeYBl7UDYuPXqU0T5NHc7y3HF+58pP8
9QfWjRGHm4PUPOIpgA3/3qCMg3bk5V7TWecL8TOzv4fJSK/MEy+0+bcHRTF13AT1PmkB5rDMqDp5
+mtD6s3SmJdtqDLC/sG45BSJFCcF3Flf71Chf04kkXve5ND1vrUNIjQm9L52HpyuK6Tx153zvdit
5VXXjpK61wnSknmMeSHeJ7Sw5xseh/bhlw784gBAbu3DvB5Ei1Tklv38l5QuxxfCyFH6ViaJl6+3
VaILDZJR6v58qTYUfbBmApaqI+cEKM0pdjVHncSofhOxrY1d8047gtnoVKkzua1mE5jmNtOOC53m
0aw0YdhU3DrkQatN0cBZ4C6bvgjzZjD6cBrCSbHe8PG8lMK0L2aEFb5qnzmYITn6rWJKt9Gy3UAu
59qUxFEzWu8GgSMPAu/eQ+SAcsKYietoUi3g0MlHpoInJGVSsypxs2/bqH1opnYdh/fzwb89aiSW
qgCTsxn5KUvdcU/AG0xFXT0hIYFZ4t66v1SQpWTnPhI/vhrvLG8k3YIZqAlZ82nixtejHH6elj2C
Bj6tkrSTbSOlUZ2tFSaJmhEd2zG0osAx8cvCdwYycqhKnQd9rwVAKOvbQQPvS51DPs9uiBfQSxyw
hPrMgPL6drbVLjg+VeuFq8H7+GIixDh+N0TSaCjOhJZCn1xGwyYEqXRO9fIcF1pXaAwu4wLYWajp
NofuBwZVp1qrhdUQZUxogsfX6g5WkdP8oGEGSwkidMzZKvTfwgEV+TIMW136kutheZ+ocScRmrjx
8fkje5+Po8OSxIOoPGQGeDXPuIoqAa4RUXPrkMs4a7bhRDNw3uXTYKVdG48B5ruZR1hr/ZCHgMMq
q7RjE7l8jWznZ1zq/CsaJfqXbOHlI7K3EE7lnjfwBRrc5o68jmop/pXueOYAyirf8jeVta8s179b
G7bXATe0DCcfByARd5RNwe+wfg+kIoLzb17OKxLFUKyOTrVGWjTzhCykla3a2XbaBnagdYf7HHQi
Wd6lhHJZmBRDwPlP/FFBMfmj5OnOAgSJ0rahnCotPRMyPAjzQNWwbMjsnPpXzYArg/ZIIJ40glwc
cNNvrq+GWOZlfF29QdQPj4ZRnl1LMQK4hUDjjMGt7V61QHefSvEyJyzAdsRZyxM71mzraXbHNxsA
c3/hqFF2FYldiF/1Fe5XPetdXfZJXQn2mZmO0wWdXq/sDcMdl3yO3z/edLvvFtfQCi3BJjxUHFjn
1IgRhC7H3QSCvKwCag7xyerv7VPfDLv2FlaY71Xsky37je3OdUqxaH4sD+kpEqU1fKJjWYoUbe3R
xoRX/+ptqfy0TObQCsYqSjG+f/+HquleM5n8h1QFDf46hOCvmDyc16oza6RWJqaHw8ye8yGJSqLE
h0m4Kqdl19T0NRvYWfpvFMg0aCGtY5dQ4lFRMdGtpDk7Bo7+kjD84QA7vX/mlrqIOBPtIlX8mYeD
RAJ+eq7cTzwHA+Qj5ilMIE6fKY8VVB0YXC34PZkwcLnoT/+xdphWSNqT3/fr8muFyOWDi/WgpTlF
S9Lil05+OSj5j+lfmqBMRLucRbWC+FBnQRhhovx9YTCs4o97/Ph0MRzAb6HfgRtC9xNK14h00ZRT
CY76rl7MieToIE/A5q6MqRGrg+zj8E7gMAlPRgKQvK8tCs49zi30vpfn+O1k1srVB0J90OEiGy+j
JBvcVke8DKojfCCd36eh3abc+C/reSu9stX3MRBfa0tXyczWs8C4PPpZM7slhCg1Em5PfPulUjXW
RHudP406RVC99lNTsGZa9QZIcTExOJ6xIIzmw/zavCo1v5msUGCWKQGbwSZJ5ZEOnEuWBtxnORyV
71eCvmFmoDYvz67yEhXVDyiNkSAbVNwriaTwz3QffQsqrkx+15ZirDESD18tC83rwR5L2qZc4HEg
UYhsSMSEaohY26jSYaQeOZjBmp4lUv2JjEBDMcgmlEGyPh8+bvYU9PjMaXbd+JFJB9va9OzmFRjz
PdL1rzn2vRUaNF8mRtRRWNpaaX7Du9YKsbnao25MluhKIjxpQ0haTvv9lOy2forA8trDMcXqZWlC
aXMM1EgYl4irZwYlHRBr8fEZLIE3SANu4rqAWpQlo1UPvrAyYmC/l57URqzuTiEpAxUYPYe9ZaqW
Nz+tLWLQ5VLrtmO025ZdNHvOyAX6V4uGghNEPPxVG7i2pJ2WZ0oUQySgpRb18mCCgz4Z5p0GmWx0
Oa2khlYSkugT98UMu3k1l//X9nAdvYplGSisgHBJoVVBJm1A35Y5oDOiRYsfopaalz05U4k5FYul
cQpit8ZwzMrWuielujnlDWxUz6lhp7Gf/PUKXCOv+f9FfQkCM3XKmvnkkbnMFYSAvkhhcZ8NDSbR
CciNWYD+p3tsw87EDRhsSuOVl4nsIgP89xuN+yHUry79xu1g+39HEdjY1KNTwY9fu8rNF/vf40MY
0lJ/oJoCpK93lpQeXA8QYuid61qUng+LFMibPQyDL41LMh6xXUiciNvvU9CyCPLaGaJWqYf/6MG6
thPDGtHlARBPawTSTKcfST7T4KzHUm4qq2/w+qd4paB3Xt6Pp0X3lKIoFruMDv+JHaFwk5ZWXZkw
joT9ylECKlwFY2aq0+lDQ8npJnLZn+Cjq6lKdGO5rDvPdq2DGd2MyYspta81i2i/nUKuzWV+DHGP
DzG/Ux/AKau5SniuMoP7kIQ3v102lLXMVjC3MX9/7GH0DtWop2t2ki9p0pnlszvgPYdLohprQehZ
QfIXpF/AU1dF9Th9mfsxXBXYa8C/qtQIFw9+l/uztt8UkZ8GERHC9gsUvu3dXs+nkPia1rVB6tIf
szYN6Z30boigfkY6f893m7uCDy+pnbPwCz/ZKHVf+hDoNGQgBTPY1c1gfZR8H3saO6OVhEd9EyJ0
Hlmt7R94A5nCGQtGR5t7pB3DOjbNv86t//co5V0FZApv/myILfXaK83pLSKTfS98yfhQWTHmXU1s
4S2jb6BWUWoIWMqpnoqATOMaxKXBGBFxLVm1IeW9YWnfX3tvEtymnBbIEG+F6qZBxD/jhhOv0Q3f
LH0EUmnV/5UGQH3zKHY7GvJqW86YXX47nv/WY1q6Am8OXL6eE+PAtW5o6ejQvJffodstJ19u0xUZ
p0rZaTWRJMJNfRa7dLqtTMa4KU20Oytl1MnNmYAJPF443cOCuf8AeO34MCnd7AUdoNL0w6+/fncL
yQxR+Y5tmqpokbuI6Aqc4NwJd/uGCo4iDnkCtbVT3vHA/Kk5IKtyp8QyIWOi9+uC9yDwK/D1YMjF
fESsgp81hnoWlRp6+mUTqW+5o8I2c0EHiK6Bl/1a+BGAz3RaG3Lyu2Q/7k2136kO6/c7NB07Ap6/
yTf3jkFE4ioi1UX4yzsnCYOtGTTrOquv4Bq3wFMc0npPFV7Rnh2/h9nzAGRcAnf6/5mALJjMjlTZ
+uGyfMNmK+Iu3M1ialssUn8vrcb4sFq6Ml05l/9GQpeGSQrEjW1c7AOWVd1oS/y9cYjvy+aR9YCr
TXG50fEm9BSPzqcO5P7cNBNTU8hApSf7un6kCaqZN2vz1b8upGl7adj5Kv2AKVeexig/oGWEc1Gg
gNESIFAEi0M8t3ycmLNmmIf3QzPSW6xOdWRMmGHkO4I0Wi81T7XbZ08nP4xhzmAc1WKr8mT6qraT
AxydPHNY3xAjD/lgbc5MkOnwngQXdidglN8noAhl1L4u6353imPdSTtYO6rZxQfwlUh+3UFehwIS
b+Nkptgu55le2Bncto8mPBJomSR7qACExoOIbbSKYS7nRNSHTH99FTS8KRQKRHSVchw5cIIMTMiF
4jN3W1u99Mot32Tetzqmgbm2z5WZzgsjFJOb8c8Vi/FIauMOAMC5ZZuTjge+ympR7CdWIK4yREIt
U7w/HZhpzRfVMDYpHfxoN8HoOw66tnn8VYsMlMO1NnyN+u/lgnBTrYgriNSsWDFrHovs8QdzQ+2F
8dpCzVfQwR63FtdKqwcW6MYNmwmwNV5TiB7lLqbMTOeD+3c7HXSLF2UV2brtL8Nn1jJTaE60vaI9
fGCGFM6+6o3xRidUSaGSsVSjnoKhLu7ABTRMwTIGq25Mh2DQfNzdFLFABtXuk9awvDNvXaqZneuV
eLexWdI2H8yV1r+IWiiaz1iQKL0qomUQF7vZAV7cdjOBRvh2CHhopmtuYcbzj/x+TTuEgwRoCa1C
I54DEZDh+VeJBa2UzjusoTuBAp8lbPTSHE9eyqtPM1QBLyGix+F6WBgBqs+EJguu95VvfkqxDrz/
7H/Gbee0yJHJIQFFasjcA07YSHfywgGL+SuvLfcZ1pJt0jkfG6NhYQr2aThVQY8idnw1Fujq/MJc
/iYWzQy3RV70hh6Htz0UJwkCXivUVTcD1V0FRRgocnPWAac/zoUd0nFhELVYuHRtDtSEYa15shr1
tEHHAQY8nzFLuLCMbC6JBs8kM5SX6nEvVDwLaJP9tM+3dWWz+Ybem/2r8xsPrLoOahztw+bV761T
JbiO4YSbBoWo12/17giQMfH1HZc+Jy7VWMeVHJAtyyoHWA4c1a9XmjnmQ+3VY1oyS4dDjOVTvy1U
qIhjmAN5+dY0fBihns5QJqABpdWv4ixya7I+7n6l5KQ4R7rzoofWgwGic/NxZqwnMm74x0FAJ9aO
zYPOkEcUM5+JrXMba86jk+X5VhS2/i4CHO4ZBN4L1qjodP+Hg3PigCPlLO/LlvSacWFI4V/+IlwO
aLe/YLNDPVMoW0+Yb2lIccLNLYpUc5bskNVWZ/VNt+vjCtntciVO8FBaL4PBoXLTsClfbYTVMfiR
5mpHlDbn+kunZND6/aPDUAUrf1YMSw7yb8LF+X7i8oarmHQeqnrhA3MGFBUkY7Ia7YbJvgS6qmmL
xNLS1OjsbTkCDsV4gRB+innlE8IY1ZmpCTodB8eF2upfUZH3POuTJIzY9aruTI7MPWtl+pQefEc1
7/jWUnALXF5JyfxuwnwgEUrBEDAax7kEfAeW8kGQCrmFCm/+ycLoDLaFB5hDzrF9R1DCj+HYYV+W
8jEIrB2B4ExdQjf5FPR9X4AWVQ/4XQ7L1PtUnvqOnpgDGTBsU1jbwtaGXelpMqN0FW6BYJL9p768
hVM8wpdodcxElzxbbTWNPW/7TGHXt5jEW0dcA2FzL8CCr3CR9Lj1h71syERJQOLMz9mbJR06WQFW
m8p9rWj6L6L2EbcduJkpShxW/Xcq7vkYi6+QHvlx47No3CweaRxga5yTaePlR+HgUTYb9Js+xW7o
+llI1l+7zEy60BDuwAj2deauXwGi+AdaayqaYoJALlQp0sRsEwNOG8XqkEi4L5cl0tZbffbLVPDd
07ZODFCMEk8P9MHWEAOjC/jkw9wygAVFrC1p0jXVv1YouGJ0SNnqLWYBkwaqgFm8N5tPYC8KiCRh
8pIHv0bYza6UHXVTB3vDw+b2sUidQX9m3WqKKHU+wZPm77DJSlFdsnmvCN5z5enLqL+/YEjflEd0
DxlMLC4OFgDIz9Fnw78+Qm2B/1v05cVGCffr6zY3YuVJarz4AP6F0ybebKotsTNrhKxvk8crNeJy
3yj31EDngV2o4pMhf5vwJDx060JroE6vm3RrGPtOgwYd435wSe9PHXn7FrEMIp2O73dDhXHzLgAa
2DFKn65Wy7oMIDyFkqeIwAaeZL3TFCRQc1TJ6UxxOSnDVQkxGXFCHPWV+UNiEg1KvA6y3gDNSQi6
BcCJiUQGtj3sBoJx50JGW1yc9jDHSCrVQFCCfE5vlGZg9GyXTkBSr+TUwC/pEXaLwaVHBT9Vpji3
5trKYwLvCT2wIF0erz/COuX184TtoIZsc9Tx2ktyzl77Ll5WiLU+/Gc2oiYGjJ23erRIoMrsNiht
OJXH3Dtk/kpedB0Gfq7c9U0jnj3eAEPiJ7ozlXIZwlODZT5/pv3S4MVQbGiPoYXIT/9nPle4cJkm
QjTP5GKnVZPGmu8UleYLe2FR+nJv9Ney7MmYsaz0Pxt+1aOhfHW3AzZuTC5Ov0as+RJ2jfeu9lQX
YNHfHBpyBrX+m2AZwrPuG6i3J1E3pJLdJlvrCMkqumeX+EUm2bfQQW35Mby1Km5UBexxovEBa/Jj
eGe2/ViM5XVnJG/w9CiEymY2SxuHuCwCLXsU6RwwEBHygMfJ3ZYAlgyLxrBo5glipSCKdduDpNx3
WEOVnNm8M+8SF4f0ZtaJp1oAvynNyDtdWPGstzPIKr/RmHrhMnUnMX5l7LrnPzmnx6G3zKL5lT1m
urjv121VOMqGDpg3qL2i6CsYlxJIyPULkUVyhP4fVvFQR82QjeJWwkOqLIfQcUKtgoFxdL845vWg
QVVBHyMzdAJnDMTyXKw3kWGMdB0fuV9gFCPwu+v+PBAyDBMf3GyY3waksvLjp8prnJFoSBcgRYww
c2RsMue6tTGTWWZKqKjFsoDzitJ8pat96xjOqm6bSOfXxiqHPOwO9yPU4Z2jWqdbwtQvi69eZ4B/
3bJEIRCqmlE/f2BLvfjJIVLgbDA7SdxkgR32QhtjIGdGJn16HjcKkUb9H088/y0s8jLPv6QMGkRX
O0ackPs+u8r16VOSxj3dgPajMo+kWnYTwLB6dyeq+yYL1UqmhWTyP6sNVi5aG7Zi5gn3mLTJc/Cj
1YDcii56g1oX1lF5TRgfeJcezgT5slrc/B47lGXzsQz3m08dtHu0mcglMNjnBjXRgaVgZplbGyBj
lU+TNty+i19ZGucDK3zACHB/0CWf4eZFiNas0XuXUYWLSrUy/LumlJTph7ZU8DlwbEHAFf/+WjOG
El70z0KzCU0/H8fY78AfwjovfjW4TvICu0TLF7T3++v3Ld3MXwes/excdHdKERjdHx9k3YWYWUNp
7ZfX3oVPxl18n3tZPW1EyamNUiJ8JR+j5svLB8UIm0FwLC1Y6LlLgAdGCwBNDa7mta1bWKLNG0cC
pmc7l1K43sDIz47RCYp+lyIxv4epLWR01v0f135zXGaJUPobqs/eK7GwgMcJ8LsHCXJ7eh1zNNpX
IfuuyGf4Fa7ZlRIEbZeB/QyfNZZBAmiEcQG8pqyjxyDxL7ocspR3pAQuKs1RugulvbibBNzc5zf2
ZX3fKocLtPajHpH3P29nO4462PxNbEAn8aBMji49Z0sxCPzBlvZtYLGz9qjUeCEKVkRfOewXmBK2
s2O3wsPOyWA3eJONNvEIQa5bMYSiYd0S1dRPUPcZ8tTQ6NFdX6BIj0UtIxDFb+1UC/z/UmlviFj5
F5JqeBq4d2GK4ICSyLi65IU+YmWxSrzO0+nClB0oSwQ9gt41wq28wpq2eP2Iddi2YkABE3edgmyo
9Dt6/XAeUcwrlrNID6RoeWIEoOpVXJB2CoIMwRDd/PcBmTIO+WNK6w2LuTLP05fxdb3d7FZLk+vj
yCTXmBMEOQ67jKLckjxldHbsUbRFq1ZB/9W265muKISiSVT/qINFXwHpCRnRW7/NMHHaNKYFXJZt
8/ffmTnGJ54EgbtJIyBU6Rf/b7HIbd9lXZ1xpmpWcEmv/ii7nHpxiKUZ8kdH4an+Tm1RIj7cbDp0
Li1h0WYi2cE3KwVOIKy/tgGhdxlpT8E6r2f3kKoSLlP4MPibptfUoyRtJYQiuJvwWHCVRBGTSO4C
2XbBL0qUkCfcKIgZ1EidzpOr0stvwclfm6mmtFxJZXmB+qZJvVsZXDD4HlhwXJqY0icV102M/e4W
0Kg1QOhwP5nmPfnmiJ3r8LK2DdUknsuVWSywinacxytxPg83Y5yCzqvK+3KRVZp/+O4vVk9ZgXuv
2r+f9JT47cUNIOeyLoSavcEstPcLAGaoA7zedjFBlipeslPnwHudStkqviaQeo+x4PLHOfKb/Ezp
fG6P2f7SBJ0S+qO8PQkJ49K0AeHLwTP2XezQxJ+yrY2uQlPshjPvd/01RaX0+ZaSQ/JEYdW50XYZ
9kndmiUDqB1zOK4AAmh+bQY4BJ8TuCqIFhnbhB+GgrBIcnyPamcVZ1VkuN1jAnkyJHcd6c51nXhQ
f0akslI+ZqlYgoPu+e1qYeEmurj+YYH9bjsfad0sjP/WYNzXVFCsHvUJJz4XYcRrxbRcfhgs4aWa
Hq98Q9239Mwnw7GRuNlTIWkz+XGEShHwg+Cwjnw77ZlzXdt4pJnUrC/rCVkEZ+/ktc8PCqc1vHHk
93ea1quo8HrgcuWRWoSqChGl5NnCbR+ox/u+HP65mzh0X1FHVSR7N52z4QUyroU8KU6XZsV2NYnn
VTu5sUiXzFK3/NkgBmtFCukh1l9nyBy007e0BZsQ8gJgj61H3Rpxs48RfDVmmTErk/TE+M/cJI6V
iYO7CUgwhnDAVa41L8bbCDyWwjmC/T8MWEgQT56I2yLU2pRVI4c8Ug6yB+OYsBnnxkz2TsFag2FP
NPmI5Y/BhCQElJTQoMx484V86DXpGRJurZyYuKxwQ8v0rWTdGSBuRggWzFBxVEoohBxuu7Ys72JC
2gR5B01bzeqR2WXUKA1R/+gwBww5TGXc4zjMuCmXTJ8GGnHpTLfWRToN5bOCoaAUmgw7vurSb7kp
BYClCqViMgYNNg/fhlXPSUDaDxFZMYLIB8tU4jdq2OsNxYV/fm/yLiOC04fJ98+R5q/h0gilrUGu
1cCNTmlzcphuMYhWUOBAeEG5Tuxjncw99yOpXp2tsvpYcqfWJ24DU0vYlcma+MwhHhDuPPNIbRXD
UBUaM8Rxq8VEI2K4nbM6PnUWkI2Up6Iqhv22aPKYlY0jBHj2pg3/NzW7N+wUy6MaL1TuA/ql/EXl
SKWphhlRQcyGX7Ef6iMt5mXgqoZmzctVNW7RvsMRs/963ZmCZPKnLr31BGuRH6jYRtWcvJpJOUDA
lYzHlj5Ls0A1HWou//dnCN+I344e9Bk9hzAtomBozdK5SLK5KRRw7myPBL/nMJ9dzzgOTTE7YpNb
8syIcXFjbj4LPl7lvTd7OSfXKcnnH2uCmKfJHTC/JBI0NFUf0rpu3R+uMoslmR3DY2o4YAfvj8vE
KBNgJazrZugSPqjR3wZ95gk+ThRYR0wXmhZTeJhe76UnLDgTz4xI9G6Jtxs8+NVsH8zLsflQ9jJm
cL58W9zK3TGACjeEsSkD23C5afGzJEO/jfnpS9JrlwOtVETWrIwQMQSwE2T16rTgpVrnSxER7ByC
F+zh5U4hZBQFODYkaHKrcRxLoTGG5uy4XAsrtnpR7iWBsLNpwzfpQpKCBRv2oFBFD9ipabvpy3xi
T7nhAMV/Qdv9uWa9qxVpSSYvGiUWAMPRhHrfln1aeV//2V/0v92vTO/sDsG91ALQNrxn3nQhJ9J7
FVQQQg47jyEE5t59oHAupPNZ71wfp8yOjUG9L4UtUxHLaUlpiW9w9pXJPBEKZf7XNoPRuPf3Rqe7
X3FyKk5F1xu9S+2lDJEwu03jN9rS3urEi5fQyWGZDY2z9xfZe70ZJ8878PdWnYsfU6E24Rmq9UOf
1UqjW+RU5/OwPtwd6JZyjsYdrXgfUdWjcBqkPYNq2irSxiLPuWrmTlclBYpXFsf1mNErOtkb4YkC
F//p6Gq5cLc2OzxeLmubE+2sL8ONDqdkV708n3TpYADL+2EawHz8O1uVDbQKuFffbhHes0xzvTLP
eU3dgFiQ6qnwXuxIKEuoKf5HXNROEeCKkhq6rodc97SwQslff9iP3SgsnyntirEqXzci1k80eSks
/Ay8Mep6e5WsvbjAK5bdfTNhoypU8tEaqI72FtRZghYtXiteHYXApG7ZDyva2JsQP8UO8QurgPqd
gk3FCefsUWTWlsbVEVcrR4s0bUvGeqkuduzhqXhoAUz646hk4PIkwJfqpqE6PJZaC+lxTGBLBEdh
WNUTWSFcESr81IjtjNc7KBw4LPYfBGV/To13mwf8jA5GF97EC5rC3B5a8oL/Kro3pEk2JZiMhwUm
PEbn9hDX/TGWDeKaNegD+XsHiKMt7O5Z28TADiEeVMObOJbSziG5bewaxWVnknx3BPxUlbOtoIF0
VFXNMRlqtotTzZJtAbUhham+I1JLQ31UDZ+9mtVn1oo1fjl8RZLh/N37GCyd1rdTcNky4Whibs1W
KyxEaiBgiZkghpy/RsLKZvOT+5vb3tONtonQIm7IxQJgTTgj7Fq5vJOWoK2lVw61RasXLGp8NdeF
JKIRpMoIY1T5gSsLk3YaDxAkZEKPNIzedMNhRLLqDM6/yWXGBo7+enEpAZiUJtJnotW9PizNuc89
I7VnHhv2QDzMNB/YjCw1tZNCW0EdzJlcKHg7cRxjMPfFTBF23QwAvA2k06057Gtj4jzMjzWUnHMj
ITM2Fhu54cFFrZ0pQo84p464SIW3lOfl20g7sq9U+VUlN0Dcwl+Vc9UWzZwaZYaMpIM+pUVFhpHZ
ql+Q5ZFDSV4ufa/b9SN6Bq17GxiwwAT9GIgN6EqKNd9oE+xiYWM5FdtZMSLLTi7ynbpcUZaNuccg
99DZpHsUOCqnhLNjJ0c37mUuzz59n0Al+OC9u4tgccFSGYz1YCvnYuyF7IuSOqwiRP4vlhW0durH
bLs8YndbhqiXPAjEzDm1+S4dch2CzAvHZC27pn6ki/YDgd5cOAhRAgiZxOdJOulJvaeaUbOQAJ5B
TBNaXbjicvqVGZZCFGAbhJPJm5bzUofbMUmbVmz5e4IRErGYdXFp+K6I7LiL6ocrwd5pRxxq3Gxz
tsPIlsdZcXIO+mmG+ODjPMuMm8bLPnwrFPwfVff5xR2LM7T9pRWqzV57mVLofUNFEESPsRAlP3fu
Yox4Zzm503VuhfzyVAa+CKDEfUeSV12eRhGM0V4Duo2v0SzMs9n/FM6SC+VzH5lK+k7g/CRqyVRx
/jbji0eP9TUBAtcO9MgAzrfSCgG2JCx0AmCe3CGS8pNeQRWWtO7LbYIrsEvkXKzgiNQtKQOSnIkU
u8By2EuboR41SH29Bt/V9LrTvxK0JHzb01uUHOqo3lsqLI3QUSZQqzNSwuXn0ioW0f3R+ZOEsGo5
yzFMXtx6oUTl3XEvD5GWV6LT8UPZUdXk6MHt3aM0uZLpO5v/XDemr/SDtb5CV16/a8FD8MYtz5Zz
yx0pstGyTwgu75FLmY1Oxmcj4HSNwgVKSg47/Lec8OdC5lPfwrAO77dEFA2cBft5/f3I7BqW3934
yQ313QU8nhqLjB79a9fgheM70j9yGSpftDqCBokbOLW2Twp0LwUQew/3w8sEPhPh5xH4vDGYvc48
h6lNaRE560Yhy+qah3vSQs6mFf7I6s0dJbQW3tPOmRov6ldMV9xYenA5p43UKbYLETpo6zp9ZW2Y
DuIg6evyr0r7tbrOBiiV8ftXqNvAMzp4osC+4xfjjmVapUcKKI5NEX50P10fLdqldQE8zMf0GySn
UO5X+DwxX8XbprgH6Gj6pPP38Rjk2cdaqW9IHyQ2txEEt+O3aorhzD3TCZXKGOM7gJNO9bKlnP5U
qUdqTI1/trWLIGnW7+nmni1/Z+8HhATMSdtl6IUZBETKoFreBomA+nz0LS+NOZapfoDdQv0Zt6eP
vQLPI5nkd0P9a/NGaori6IqMYITVq/idt0TOwlwV/IuFvTN/Vtyng3ffQYeMPV0tsyO5UjFVVBU+
8mY+b2Vty6sq2j2S/AkgfhRzv1KFC3kc/WfeGr8in0vKOm4Ox8NBQ5ZArWsD1T7Pps/SPooaU/U6
zuOsU4i3RrZd0PHZGYBmjRfIbIGmVNx/x7iAp5sKwCNdjwMA9plqqnOvE8lKQZvpn3u7uz9T0Djb
ilX3oCXIoItttTP0ZRimC5kGMjZzSBw0OLcvLcrCC+G6wyyj6ePs4mLzP5M4cAoySImEfeH3qjbz
mSyVUZE2J2pZnEDbiuy1s3douJQ1PBRYEBs3RUU1lbV3G0TL+xOTgzz9z274kQkotI+oO6+Z89JI
FOUYn2spHmpU/9Saj6sTwFWhcb90B10TAvp9bDupEl9atN/FEkDFTuwVTMgNN8XwJkWi3DDXewFW
PgWhJG52gkIDb0Kv64QI1mtXlSo173/1MDCvGpy7Khfs0V1/lf6SklpVvLPrFWfespN7hUwLlIJ0
tDVw4CvWTQBu8aj78UQs3WbRlfzVVfzz3jrYDlULlq5bkC2xBdbBWm4okx35QgMVL2bFh8QugXIu
bxN9VT2NXGl1xBMWM5ZUoOmxJrX6Y2ZFNPn7RMCUhJHY2fGCmgViwsq4Xg3Wr+BvitB6a1aySTlz
K8BOK9qzH2dPoLoui+urPI3tPvY5sq7lIN/eBaIyipVkeMxoJIL8W0SnBgESjbFTbrMQMalQeXQV
bdChLF4w/2JUW55jrRBhJ9t/4FClMefTmzoW3qLcU5GLabx2+3POgoltfvRzr3p6pLQOxDlwKm9e
4ybea3dlQCb8fKIW91lyWvtLvxHWhlnqdSAYzFSLIP44FRggtBAyPXYFP0rcGvP2jd7RAUbukyb9
42dY2BNeqsDEYXQmAKa8oSZscq1lyx/wRgBTihf3EQRiidatnJM/CNLG295b9P/xoqwgQ5Md9dnq
2LCSk+SmYg3ekb74fUOglABppi9/ojRAUy0nq5a8KA+0eMeIxohjHMltC6KyCvZGV8h1l35C7Ql6
5CD0XHSm1kPQDPxx9L8td9ECgqEgjbmzW8SbIHOUszRNJkv4DQTGKUmSVqVdWsOGsoIdeHgmZIqX
VGNPHO8CeLN1QxUkx1XJ66ttRW4JAdRK9ZzoVUjEoYa5Z9KWvBkzSXQg/sAOMvsk++3I7XYFiVKA
KosWHliA69qkKJmC0DYUGRpVJveY/a9zVgsi0trKGdHLr4h/+Dbsw3MkZPkg5a8VCIInCYfe/yql
sLyq42uYp6JDcDlfm3JznuCcBWOolpW3WpCzQC1Cqs4coNB93e/M+QkWyewUD2MhyeapfH4YrlwB
eVoC+N5irV85II2RH+k86d9qT2Zlg4gwEi43Cd2a8pie/CEv+/TkwIeyojCT3a2K0gb4N9Wxbcp7
NKaOJFWOve07qN3//W+VoDmaGmDMOmKoRMqoPrZvSEs0Mau4Zv2bFOIcZ9yAyPPc52ltq3lRZQlc
Vq7gLB/gBhCIT/0qG5HkbAcHW/nvOdZZcETlnRkrJtylOv9u5w3KPvU/SYKw4++gIqycS7trSD9z
ikJBB2JP3vMtcekPqeRCOhEhTghQYqCOLBbJ0KcpySTkOHP7RZkEa4vH9z6tp3eb3aWfj3vKKh1X
t+OStPcorQ+Pyr3WOPXXqNmu3fBXYSb++KJ8kvmvLTUrYU0t6l3qZfc9MTwjrNsfPw3T1v6qgo6n
o27YOciPd5rqXbFK0r0HhfKywcgR9NvdysVvbge7LYRwkiIWf02qXLlf/dKTMEHy7bnKRvEzVuje
n1oWDaVu4dLfTuKsvM1/FcKHMTXmFkGWfS513DfPfuUg+RjdUllYiu+iHNEIWvzWNPB/2CiQhOrc
+hmxYd1XQCo99E/Si3GRWvi/bRtiBgj88ISDRx/4O/Uzc8kSHA5uHw8fpD1GDL9c112ukhNoHaLS
dpawEGx/f5S5PvinHk1erfNcDsrD2+/LICTEC1buFXGjSbYlPnOMs8d2de+a7yrePYECD2kryXc0
B4lSb+T/4rK59XVCeq9nwv9rULdSOBVjGM/JchmJbsssNv6cRPgeTSlh6HU7eQrJf1xo0yOK05kl
Qo2dlK7b7i8DMe2H32TkYoMjkX4ifFKGXx1jhp00OEfAYz8SGn0KlFFKoaXmfJ1XMZtp6ShFVZka
IqHcEm0szYijCNuqglreCWp7FjCtXzJzVgKPAFNXwHC9YwgsNcvl18h/cUZBe59aqK5ZyHsRWp8F
m0Z2Ta40KAyYy1jhSzH/lx2X9hsuEl4bVaeZE6gib2DbBcALxc7lHVSb0SuMkjkbXMAFi6WMItxa
csVwV2UqoD1YoBUP+wkeSGxjiKU/+OnEZMQjWVS8zHk9Y8b5u5Iz9pjYqT9/myP8OLuyiQmfFt1h
Okw5MvshDS/hMmFXs4C1xNI13CZFr6TfiqquOC4wH7awuyLPkXwF0i5I8K0hcKMYCt1WQqyrdkF/
C4pQmQAehjoJeIxy99XvbAYLi94ifl+dm+gU6YvUJuUZjg5Sdou7lDJvkkFDHPQc8cmqg5o/As4y
6yhz8+cXMyPMuJ74xUSxLcQlNjG8IPNBAYONtsPtvqAwdiIm7vw8JFoQvCkooCpQNHO3l+oxkAEn
PLuklpm1x8OqCETMZjTl9aRc/EaPf/QadhnP138lkAxGJDoQRb3wy6jcR4PYLfEfS/4oh0h/HuUa
oKWaulW4QGtr6IUgvzDf4/IoIM2HzxMGeOoUQvzErnn/NeNJmXn9dfCzVMniV4SrLrnhY+LQ8bms
XAlfQ7abQk3XUd9hXJKjMtcg+z+AEjI2xuG+PTVfNG9Lam/pEWdbmdMGLT93lxajTWz+T6In4vKd
e2I6poOchsxRScK5uD/EoU83WfLFv1KEIW0yvh4CeUDpUsIqrqanF9EGiO5rwxXf5GBNn3z63J7h
jhEHFgUuR4TPk9gbmNq4Un2DILq63Y3xtHMxw7G6ieL0DZ3qADYq+fLOBJPT1KKuZPWP5JANiYBQ
tBvlCKrF8lzWrZLfwyRtaaums6hKWk9R7d0NQiFIt4U2GoiDbOMMWfQGZa5nvk6K/6kIsx+/7Dj5
DO/ybvgVvXwyMuZimUWVWdjFVa1zDPsQGccN3a+cSciNOOZztZD+70CyDDQLikLuU1f8MRXIlG6X
29yInHnuTdPpls54ADqdtzcrKhiGVdrrhQfWBy9AYP7J7JfoqpsBijxqOpqwQnhqkc5ML2Hu4Xxi
DDacc3U70jwl82FPJ+J/rq0Y3gfVLBnycnFkKt3foP007iCRDMVL59iZc8fNY6mORlcZYopoSNaM
dcLkBzVLDMtatLpxouELC9YfHJql6QfIKR8XRCGeJQT1yBPcC9PxhaI1wFBYuY3olGQR+GMxPl5N
POQ7+vPg9abLKn2D612sWfDebTTVJhRRSKmy92qguXrBw9xYcva0iq9Xx2xVdYTK7I5hFfdIklHL
nsVDDAnJJjteMrfUFia9kJENbljEPTK6br1SOrxfMkBXrJtpyoIpUNR/1PyNeDW+gFEyq+CoDPpH
rnNoSYHe5rYWfBB1CLb030JUefVBHDzhiMk9y58obykIBctQQMirbQO527uUi54Jhti+mDkK3w8r
jssLO3/bl9MkR9GOfgcyEb1UAx+MC5LsaDXAZTVMgPpSVDQgWsvWUWwJTizStetrbGBzqGmWuIvr
/eT+eOdWjN0P4lK745s8M0baQtxIKYeTyTRbJd25v4qF4r51W4K15ptqsr6zdKNc9KdXviqcfXVs
t8gvxA1A0Tsas0OC0TSKuXTfom2I3s5wM3WZ8tt9AZUnkfFtMOM2Mt9ew6WWX22iroJB6VJMm4im
fd3zdjIcODsQPeRB01SS1NR8HH5WJr0dLnBVfAv0iQaeLPVPaIUXsdE0MbR0P5B5FaiD95j1hoky
8ZOz+xRF8Mf/4KP6xaE+yCangDVlLGSJ588v8xgK8jfhCwJu5att7VQ4igkl+fV+sNzaekes/oaQ
f9XFZ858FS7wH129trq99h4D+9THY/qWcOnkauIgMS1uHPf9CloFxapGGokZD2BgJ/reCwqxkJxi
6wWmPVoDTROX2Cs1Q1L0hzRZjK/enRId5wS+PAR3zWVd1rF5v1eJt/ZxY/t3sE+2woBMHUHDnX+s
tcMfvEmBtHWrtcZTmm8Qcqtx/Qt4HdpIEJqJw/KGQCMzl6wZZqfX5YSRxfruivEHegMjFlyMRaYs
boB6HW952UafhEhpMl6UvoAeD5OjyJ8RclYntE1mABwRrusSSlNBYtwhKVJDZ5AhkQ7i5RwpPUg5
0c1LXr16r04QXBJTtQ7b64ucc35jOUE3KvLdOwl7qfyi5K21qR25pHRfIAIpb+VHHhX3WwTm56qz
7oAP6AaE1TUOWxlbVOWlfIiRAsW4mdxWxQ43FASYr8A3EhG1Hbh+Wtl+5wP7ZfvVPNIgpD/o+dmv
H74HpcmL1lp7HDjg4Jtizh5iyfjhIr01t20g7eBYyOpUD80XGRMGS5AJb2qhaj7NKnP2HQoQdRuL
5/i0ChPHfkOqGvX//Y2T4ccGyaktYEt5qqufE4jw4znKnqxeq8MLJLP8Tt8syeQkLaUyIfT62U1x
0m7XKh8BZUIrrF7bWJoF0S5wWIod19ya4GtCJERRzAgcPQrE8oDHyluo4sI2z/9tgppcEU/fEpzj
Vph7/bA7VGlB89zW2tu7RC8QS3joqvJtafoiuP2QeUMStcE5Ob0os3ACnXicVj0HPnjcQObgva4S
6r81WHxr9chZxWAi9ZSTq7DIvdGLEbbjKCtadYbZvCcvSbp55Z6QkeJQw0GkvPIuwJ5nbcgz9S4R
dPB7OyMLs+902cp6hu/B8pA7q2PBpuyscpz4G2A+TlRL9ef3Ld78lBfxOPqvmYMB1Ip/flgzVn9/
SFFpb73qNC+dnH91R0ti6ntWiVN9sL647jOhKMuS/iK4AzUfvRfiEvjWB6H2cW4CSGjPlFftubd/
/2fnZlW9EPjnAQ2nH6Bs0H7MdltaY2Q2gEx2PFi22ub11naiWBZ289uDqXyp4py5rs1ElLRHHmB6
47PCSV5yAV2MD2WiV09PdKWg5OTGJLz/ix52gSBX/ABJim0PdXg/o+JJp4bRTvvA+3CjTe5FW5n9
QzatbLNovkhzAI288z1Nrf7FdAeOUAxQdIeD5E/59mAzNvsuo09HN3gwiDPygBORqCKWJeoCfvy1
9UYV551d5jVBhqXst6Vv+bv5rcZEh4cnI3t2yl0RQO/BTCQrDub/s/r8wWnOYoyG8eeL/pb8BGLp
HXR107MbbG4q5XB9VeHAVjeioQChIFJgdIe8Ajq8eF/+NRD91dMO+384amSrCESk/RhF++h4GF0l
976/qVAsEaWu2mTKDeXNfCHOArtX5Tl47WMtgEtzXiJMazuDnhUvmvOd/fqwsjTsz/n95ppQC5V7
5qD4+H01GMycjNdgfsIeL+rZlis1OLOBR9fvxmR+ETC67PG8fHR8cZCR2+4hI7CU6NmrOBWYTvfm
ca9pYVnvP617Pno9pXehRBZIusHuMwJPpqL9YAiDURdyOiSeoVuki1AmtibnlNmnLKX9XVjfk5ty
8MX9w6K+1UpN03x7HCY0uCjwCpMRsgU/Ai/J/zQWcNHsrsEaAO8G9f7tcRNBm/2gjW2YBbsjossG
y82ehBZhjlppZXpV7jl/UwQWzvBVjaeaLpfr45dPKYZ2O7TomxrfmUiNtYtBSyixkx0gSHPtfB6N
F49snrnnBc4YmO6ZswbT2SUl51DkzAmx+JSCqFAMfTM4hMDmioWqvBz+VosDbYvjL71CzA1pcGq0
bt2qDeBPxemyNkbII9vurQVAzrBCXw+CIfzFUUAITiuE7UJlpQxWOg7NWrNdhi4szW01eOlXFpJY
QCvEB8LnQbw2Wrg2KgwRzDLNucjCrGiJLRBjQPMAZxKw+lYkFIfRoz+cjkxQYo0K3F7d8FXlx0Jf
U7InpHrg95wtOEQf94GWFrBupMeK5RIPRbDn9RaKpSbpwu1dwVliallTVwlXibw2xSqplvlln/xn
odGFoIAGknH3d2AIuiJU+YMYzKackosDEx7NCCjHNsBmQqjP5SkzD5XLOOuPwHY5RaM0DsVZ07ej
U4W10HWNqYNe214Vhi9shO2KgqoWQZ6iluaojVSWjl+/PdkBL8Oj9LyhFqx3NStGQq55/FZmK5Ze
ulY1glaV6uXQkIfmOk7D3jziE6Uijh0eH0G3snCsiwpqcMjSbFRIcrGg/YVOT/+l+6uL7ZYlzZIn
9Ku6F5K7g5LI1/BqRm03WO4YaV/Rt/6XUahFWRrr0GfgfH6mSphKf98gBaSCh2EKBA1saPmckApN
DzRLE59OJ7SvBgRSDtnk8KaWyAxdtUMOKup6GTuHurxiG0ONhsBZaz+M0eKw87l8UIJrGUWCLnXb
P0YJ4KJ6nbfQExdnoE2x9QPTAjXOeXwSZcwcsLIjxTYZHDvCcEstsd0lbFEDSRqtD0Z2NXMszLOW
VhehTvjdY8fA/kWDY3sgNq81SEWDh62TDmXR+BHctBWhTSYeDzGpqJO2P7E8ZlQKyREsTLIbRlY5
pN9ZhIij9C5Qgnq3Jf6I2wmREhRgw4IeoFgIPJRZDXA/hxqeEWH4+mJp3rpdmMFN2ENL/PmZCYOK
iYlMoPjHIqHoYyGm9lAm/w3q758nI8UPFWBclIxthmuwZmWAOjA8ogTDZ8nxpcKMYq8hTMk4R6sL
j9m+05DFU8wBne4Lw+KJJLs3PfBdF03Lvt84fyhktFbaWfkoAvumrGIwNOakK8ctXcmjmRjcelMT
Va0LPG3OarX5+BCrQ/BF4F23TYl/j/8yPe+oPzH3mZ/96heCmtCt+audDp3ZXtcQnLV8utBCz2c5
17HdFbXHuDX+QK0v1lLHj67ggWq6BioOTquSuAMgg2efM9YGrU21E4xb9czFAb2d5GVpz+Devf+P
nAMxllyLSGa8yaR1y0vnnqbDYNyioQzjAgU88nS+hGqRfGTKilVseAHKpVWtT6cPNi5NE8TYrGIW
8uEB1s005Xjxvegi5gQRsJZSNryZe5Rj2xUyQz1yBtuqfyfJ7Cmxc/pzt/GC2GITQpQ8Cxo4pxe4
h44qNXvbf+UBCgnmWoUhgjPWOcoLAr/703vDWTB68xnRh2tDt63w72/w40qXM17MAhXFCv9lmD1Q
TELPT2wFbQxSGHEyw32YSRXQXpVYEyVLjcTsxZGf8kmcPbynuY1umAcX51n4JndMKKtgO5j2Zwlr
c+eufFXB62uAkxM2chtuZSJZUx++kqQhkQ/PmVVJQZUUghBWQAWCs0JcRzMVbPenH0/cNB7FrRLy
xZz18xLTA0Ko/wK+GFGR6i3ID74uPDl6M47ZrxSI/ORne3Xunp+RxyG8tD1pCxrQc3WdhUbC+mnU
3TsTL+ch3WiS1OJGSg0AagwcKbMLqomjYXqHl0ey1TR2MoCXO5bsdNoQ4XkrUGlD0LwNzuBKDxP5
gW12wLxysCYC6dUR9F1ra0OCFCnyduJ2Euu93bZLp+rZ7ohtAC8A4P1MMoxHQQukA8+2jZ+IluaV
e8Tx+qyyqM0i3v/DjEIxb0yPjGPUpF+tozwsv8u0VpWaiC7AD8nMJpy5/ojnyh5gohpFyn2lkxQ1
IqQ9ic72LHofJOct92eCoWfHZhiRb4TiWFlRV6kp6WEO5fp1IToO7Px7SsWQ7I08TBoutY7mY+CN
MKdyuA+92bIyazN5WSBsaPufH8scV1jEg7DRynnWxlI+f5D/CEldxIx2W2z4PJfLUSjcoedFHYLv
tZBiw/vxFvLjvyxrByyUWiE19wbkbr16GLJ3RGTwlO/Onsznc1sO9iuGCc1KvRMnUQTPXyimaiOw
TNGOq8mOqj2uT0rT/M6hw1fb1ILB7ygghEo8fs9/ImpXblx1j5yxex9DrwLMkLk99KdR5uD8zLH/
klxtLTzHy49YIMDkBkpMxp/niwTc0tc7kvfLaXscmyey1d6nFSN4vJ594+7zHyrHFXiucEiKKU5K
nOn2ZBQ+WMe1jP4cLisrihTfvFMqZkb5+z1orgEOSUjDDhOs3wCVAAeCZklLxl8B7NRUjbAoAOt8
zsXUBJvedjciCP+2jwsvacKayVaZZtkgPFVa8nSUtqZtM9no8w124GQdJA2bE+Ali+U9XQFUIHUW
GIK1dSLLax5jzNwzfXlaL5J49PMZWaNXMoXGRuACEIlmefnoXB3Q01TmUd8+eSivJ2M63liGvu20
tkSMSZ1DJmmcvK+iPeLryr/fzMOZ+TwVUd/249/xYChkpIX/8PITyZmvL9seGuSAT9iPvL97StBf
Kt9L5xwyMEZ806iSC+bSegmqm8MAKOE/D0UjRqR4r5B3dLbpJUK4sUCMkYxU5t/ayS9EJHf7HCQq
e7owZgY1CNnjxaSNNz5Ymk2HgUDxoQUd5XuNtzgPqbupDrvp/udUfYrm0vUOoOqi0ADsdakeTmPc
ss6rYMMw7HfgfLBFvLnZwKeJbYzPi5R6Ca9T6hsjjOLETwy3duj1aOgfMJb8/8WS5kdWO4wD9m6E
FojrVflfStY02SDcJjq6Ee/KtiEdlsES85Ahf/lsLv4RPe9SKm2ntnx2qzhUXBaD3uZpWbVHVqs+
1BwhGvO3Opp7ZzoW8Xzw0rw5o4IPYTVkCLGOg7uSQZljHyM8n6jSyMuBWc44iPLq3uz5NKlAaemH
I7NQVbGM9h5S7ycQHp6hBvmIwwd8QI7BZLr74zdq6c087T5JH3DES8zauvorRP1DpIIf5ThyGZSq
SfuykXjZuZALRvO/ZSTHeDRzE1XGXeA66hD0GodT/GcuTXzcQcFrArCcra3FeP2xDkPAoUUGg0CD
RRqnS9327vkEECq2QMiL/legzS6MBynGRSw698rr+KJqYskheed3wWiGrnUY2Ne+hOyLcXh5KBK/
C1FRZ3ITgGyZpOl6QqLIm1Tz7NxaqoOneXXtuOHhkb//YrzyKLXeB4O5rOGZksOVPiWR4Q0h4u5J
otSB7q7EoqVlYoGiVPpvnmIyR06/dkTyrUhpa8jkhQxrYiN8CLL+5j0rerkUK/PCe1WkrGWNRnZQ
K36rfFzNpIErYwZ2fu4az3ik0m4m/fn89lD5SYGxqZNHyhfkTupuVu9qq2X1Fmu0XcqxdfiV4t7y
iJXz/DMz44+lu2kgYWXoc96TqNkhSys6g2qUOSsT3JG9MI8IMm/zR5njnwHVHqR80DbMEoADTEAT
uKUQqgaSp+PF2fKKl2NkEq1wzTwOCv1cSBHhv+KdmQ9WElkRupkT1eF4zvn06Ho+SH0wmYrY52vX
TXNfom+HkxK+5wAKRgrjMLkhWsoZmdknCYsmUbvhCth6FTGW9prtW9altvQQDdqDdGj/JTRPIIN/
oPjtJkEDI29oKAzpiWtXI4FxJwW1k/OdziGMf+j/TYlEiH3WgX9Cb/EYU+Iba+QhROAwAZBsLg29
9UGrYC1vURg/cYnTWDooHcRfR0kk3YX6Ref8ROyD1OCuh0iwhXPrRgd0xHRtlcLYKjpXw8C7p7SL
IxDah1j2qQmzt3siJfRKTzddMwF9tm/7+mmt+WarFfMeWaRRqUlBLMhQN1phe1GaPemCFXluVmS+
idhMOH1jS7D+CS8u1OA8B4J3PiFtdfuNCyqL8F/jeqFPzyk+jr3wiB9paEs6lddyk3nmEINIrFff
mbVZwicHseDkz8JTLoSA3w8XzHbVc7RWVHrPi9aD+Ix3z9COrXAVpSO/hzPvgm40IYfFSGjiHlA9
fTRlsYGM7HAp0Bgj2eHmUS8cXp9jpM+q+nQN5FtdiUcm2v+mKYjxde3nAIuP293+HQ/DIRadSKSw
tQH0Wptu1U1hVaevldHIQJRCKXMGc22HcHPbMkri2WNt0zQ/5yDABCsu4ss+emM14kF+gCfFViT/
tYrqgtoIM/zs3Httczjlsqbbf0k0p7N3o7PHTYK+mVR8zESvXCNIFkbGFbIK702OTQQ3m148aOde
1+Do3UFXHtMGsuBVjRNawQ8D+PWJ/LsRcvtMs6PxHfpoiomZ0J5G1B9ZwBo5fyiHjuT1TxfdhVDq
9IXYpqrmvoDfvJ1Y4MCL7TLrytbBHY5+sRYLTOuwP5FTz+STkLLVRpaDnjVyFB8bWSWjmETlkaLt
cVoaWssU0nPxo95oNBR2jSyBNZBAvncKEn3zBz0C8aiwfGRNIRtc5/wo/h2gdcVNfs3liutzRF54
cN0KnDDkkNa0QVt0BYH4Z0ifi+MvOwB/0zfubbAS4KQGya2w89GuRu3bUJIBG1rTbhkkeiXCr9eK
ky/FXaBekGtL1qOf7EIblNh9ZiOJONhMDqO7JnfF2bukwQcgjWbiW71spXRJVnoTTRu+zjST8K7w
0Dq1TOovnmfOTmZO1wzn91ahXlHKVv2WUdz3O3k3hek5nvEfl6XgbkyjkzTf2ZDFXuTlnxjncLHf
6RAAwU6jXUxuSfpCgCwy4e8MV0Ia3QIlGR4v5tpve14ySYbDq7vWbdYbOoeweZVgjvbo8D63WBkE
swZRT1rTezPnoYU1+H3JLM4wH4Ggu2uGrtaWXiLdG8eQvM1VlgxYiA6CVDPYZoqNUfZQ0RG58sio
tmIC0qj+EnlIIvXJpe2AbohrNLHl1ykCMkJwb3cRUMt85k5rYigxPD4ihsbT8i/vF+nTwz4lBmkl
hBqmcl6BRnCw1w1I/M7jl8ZWty5uMxq80kW0T8W7/e/lqdKmjVkgpxgU6VZf2KVc6zY9fbikMwwx
p41nvcH3/q3QyeDl/pXpFjS8/1/zTBmUapfK7hCMkXL4zLOCIGwKGBX+mvZLCCGjcZL5WvTD9YWX
3zgSPSaqUTA81dpJ+7tExo9hYA6eYQc68RuEq65vR8vxNYdL5Uzn9GHz8pSSxy+YV3nA7Cs/MzEM
tM+C3zFx+q17xz3N9LroWZadUm3SoI3tT7Kd3febkZ3kCnRmYx7Y+hswbpLlc3tVlDQ/VlHro3k3
tdhCJoq1HKMAbp59lyZOL4PIyoxtTBMWgjay+HuZGN+wIrP6MZZxsDjxOpCe6HybC2gcEDglMYmw
A1zxOdY+kcMdo1W0l4cYgEFE2G0Roxa2cQWLA1rx+KK8pjSiaodw9C9X2OW65dYwwQPAXseP4fnU
CtvQMatbLOMO3PgJOIc5/ZL09ilSuwRDG7EuLzCA7uvWiY4J1XvZD6JE+mtVUMjPBw1lQPark9H5
ljaPO+zbU/BmjzPK5jk/B4ErOuycMahGLYFep7Jops5YbH8px4IRkPHAcBZ8XRN4OLpv8TWkH0iC
fnMsx3eXEL4qy8xCl3JryJDTR5oLBe9nAsk4eo20tZcviTfJZfqYGnufvVWvQ/tddGNYOBX3wqXf
Wtd20o5AjXB3SOCTrLm49GBlleAy9ojh9nsHozHegG7pSHpIZ2R4yttX/j0Wooa7LYBfi9NvLF2U
0OKPAGzFn28EV0Srw0txX99LZ0veXkywV2ZO0PmlSWbgfbZB+owW3h9XeZ24pa+Fdh6IDvYIMXN0
7nJHxLw2ptPnNtfoZPo0d0a25xda8sRBXo/QG+yAPhY03wLoxzsPw7PPyaWPNgcriY/woDulbjbX
05GngSw7cXI4MzJm4D2xESTgJZgWKan6lYQvXyUVF5jewd+AHH7WkVdun93xat9WNDteHrnY34NQ
qenvFQ7B82D0cACUKmDcgrVVo0wuhnez8oPKHcU3EJxphte/nqpsrjWRWwunzbhziNuydKcpIfRv
Va8rONNcs0A8z5RzClOxUfmqhCMOBG8vprs2Q/w4M89xFCZsLNO3aD4AV0mRbsoDa+wEA0u0WJVN
RmIcWMarF1Y4zkdCKkXbs+XmUfP43Xg8Ts8MEDssmle7SdKFXgBGdNuJZT3jHLKSGKdXgxgZ0+JM
kcqctVHepINOdcTZhTe1wRJc1xegpgAZU+Eil6odtSPtY9o914+fzwq0/q3GGMlPTiXRdwdG9t+Z
cmHQ4odmQeAfIhA1NqFK5OwTbPSQzykkshEiBW+yP5JxGPyUJQdc3zFAC411SPfdh81g9OLCV9Co
5tWD4/QdohLU490vxlN6y5j+aIOn1XjgVnBqqkjCyruEJO4SdmHgbceKpgHlVUYyF+39lN2bKtlq
Om1h+02evmlx0QBFznYdl138xYvezxLxCojFZwnYN9kTClMPVlQCrVW5pqqOmjkJ8epCII7W7n1z
Azc8K1l2oQzreV35Bn5RaB73Y7QQ96zU8pJSsypuU1Uez5X6dPtH97pLGzVP6syf13JAIvsBxpGd
HJoJcqCfwPs9/6BA4XM8lIJrVC2JM8UewmLUuLv7Mh4VYYuUkBk7rdzTeVTogIYBTefF/zUMCg6i
FvYRewiLwJ7/a5MO4I3IgiNa4mvocPGZhMDSr0hWLkVsZhsiWZVGoJ5lh9Key3imA5FPSaL4wwid
f09fYLFOlEtRoxMqz7JNTlaUXufcnESnpaPmoBSLdzOLmiPA9Uofsti1WTUvqU+m97gFa/5tFO18
Xp4FqT5qc4c1SSRTwoQFmwckyfmHs3xmMibu0UlWBEBARhVFQBqm7x31tSLzSl7Ec0oOxGpD01OC
dhyDtI9zAzs1ZcTZGT9+yIuDqGOLV+XmFy8VxKLCp17UK8R2aAM/qSmyyhvY+2god/vR1F9HcrHk
BXazk7sh506l4uhz+Ekmc5LZiDdqr/I2SODEtikW8t0c5M8CSWfYJRO49XJNL/cdj7z1GQxI8YfE
kXPUffUO+7sPcvH/YNI0b9oJ5WcabslThwlPAxq0hTr9U/WQvEn6GBF4OJG8Hbldyh4XDluT4MtS
Gk/qBeVpdCbVjhfOzDZBSPYbN6nnM0gjm9U6172/9K1S9X2GQbzXkXxavzSXr8IlE/WeTUtIwHE6
tsavoHwVftevI8BJCOFGphY8pKRoIXCO6AK25VAws49NTNBpKBpGkZaWAJBQ+IP6hXnPvSihFeB/
qglJNL8Z2Gw1PypcbYgOu9TewRdGal4kF5DM6jZvy+AQncPLwgoqb0VO3QR+7RMFGmy/2Aje6/HX
H5LfsPcQk0Y1lW3WFqh4PLmaGjdW3JVes6YwMf86+0zRa+0V2x/HlXQ4EL1KNtpsGyn8khkUHUuj
TyFvCcLB9BlorCla/Bri8cdZX2L/f5CtnGJrE+OC5gmHNx+XZ3aiX+KiwU6zVw7wmdQhMp7dWoyZ
TF+1TULBbJEsyYrIpqnhTRTQJhxcXyMeW4+BY039BYAJw/AqzcQ2q7vkK/qk9L10sk0zTC7KwAow
h1RlZxVmGGGnLGCaXwcuvVgmJwvN2Ato6rJaae723fxlJ0spaaonv2x7IeflrMIN/U7TazWFY22v
Dt2LI2/4SPLqm9zGs+qMF9vDP6aa/EDrZeMVdRRhIXHlAERswFK02GFdb8fpxZp98uIvSOad1UWD
ASUvN2YMtQr/BKedC9xVN2dWj0BR7yQTcz7nU2TLCJBrNjOOXJ69hie57haGBNUCm6LDhCujBdQc
eGRwye9kJ/diu97puVerphw0hpHesdRLpw4pf7doIKLCKR9YRXz2bbxiRd/XLVeGZt/DU9++jPvf
aZKRZMgM6tmsB5awZltOnKkUS0QareE/GLbv6g2hHkbFOvb/gyecL92SLzStgb7meCpAmf/3FXOx
ti+iVP+GbtAy4bcCBJE5ruuxIJdwPaAmeQvRf8ww7tmhPxT6YtKryE4Q+gh3k0VDh87oeKvxfVvu
+0871sXYOGuvVFmhvQKf6v2XnNBaOc8X92ZtDqpiF5FxwbfRUTRfA/E7o7bYQp6Bem0qDtUnUTUM
5dw1t107hXi75VkgH1JeW/Kz96EQhYUZNtzi8XvMg1rq3IdnGW17Fyqe3r4qOEymmhTHSv9hK/7I
flbXXhvvFAdswKuEc0BGOScnU3CdIQRpJcDJPMZDn0lJO3MzNNon/mt412Pg0IkwNQgh23xX4vKf
EIGAm05CASUnqCmxyr/20k6Ql4aa9uz6w3n6qqeSuS+/pg+aFqZCXprmYRRIsVKydNYBlP4Zq2DG
inFWDikRE+St/fr4SNwuIG65Q5PqXfr4d2QJtbqwwI0dZOgbYaYmFijsi1iFx94AOwa7NCKI0T+K
xjykHxKhmDd9EEkmmu4QOpVxOzXJ7aS5KTTtVD17sdZdAsQdRlEXQWRG2DTs5Va9iyEsgJzzzuYd
onA/Sm5S5Q+JpagrE3uLDwIpSPuRPO/lTrB+6FKrxs2hu/9jIYp77t1eTOejF2VJ3UiOobf4HfNa
nXg7WAylefJpz/kwSZoVHNuL5k8I9f11TQmXu9BFbR7HeOMyws+bbX5xa9MmBivZe523Miraq1g2
17OoVtjjsQxwTfvMSkbYas27XnFngV3FjW3RVlo1Er/lnC5n4FlUadJIwzCqtO/15uAcUOY8bdWC
rSKqPibZTzRhdVMke3WknDm0LbjrU6YpWeXGs7sFHGVqJRBTkxudeZEgi0nDOw+yt+q768sbDhYw
nLgjCoP8b0WzyNvhCsGFyLNQt8NXS+3aHnm9q0gNWE6ADKao6kT4bEBO1wRYVrY72Q9Q0DO68bKm
MQugmf7//NxarzyOQ9ydyOoEFs+AdTepIGpdQNSkfBbw5ewhHDmmPAPFCXIHQek6+OLod2QSGp73
rbu54VPUavqa3Veieckm7/CysMm3HrsMOBxTzRcImBn0f7ymQgT0IlRjrcxPu1dxusuDow53MHSj
IA6mnegq/4nkjvalqsZRV/QKtD0beBgtpd7jvnb/uk+LOI/TZoOSRu2zb5xqXEwKscOMM5LkjaF/
0NlLY2WPrXHleijh9ECVtPLDbV00Nu0zRuI9xBEO/f62czxPnBLeX5zKSS23vJVRqEFRNmlQRoRi
n286ITjselWpb1aOUy2vjHvqTc3gSDPqDUq59F182HjqeP0wsCLEfGvcF9H1Dd/RMpDRYBDcdJVJ
gUNC0CosX/Ok2LG5AE3TcDFHlrNdK4PpsVRvoPNvdeooagcYkvfM4zxPQ1dB6C9klooeolNght0v
Y+2CFMwzeFIluP0gSxpYJZOwM6zBRuMwXIMs2W/ceQ3ujFhur+UhSxpuEWwNqtKw17829CUl23o+
CkRVBqYsKfHJOukBckMZB4FjC7WhgwOSlMMjX1MP5bmYM2GKpCc3xukAfQ0P2KriEMejV2WzooXR
/0B+LnQejZyNI1qelafVVYNHMVFzRoX6pIUHdujQo1jQHb8eIyS9bm3+hJe8rO4kTXkhx2SqlJDJ
nEntAc+8jh57AHyRspXMw/MZjaKQ0n+nXpZC+Apn9GuZSfV0EeLiUiTnNB6E/HuvOXThg6EUm8gr
RovZ6B+D8E04iEq6e5FyAoE7TJN294un85a/o5lPCGxmBoEEmzILUHSzTWYGc0NV2hNSno4Z7L2D
YxflI9EbtwEEs5llYSpUIJsLKYmtbgyn2iRYT0SdCp0kFPkhmWk0W/yR/97rSnA+xswnooVhyHLW
LgA04cbOrAjxdxTf2MCqj6MTENMpkrzcHcE45csJG3Kqpb8qhzgUQUu5rPhkLPzPglgjmHJnHFSs
EnM+pwehsV2X5ErJCZoTor4ah78i8CaosXMHuF0OhdwRORCgE1d39RJNvc1zUQI4qriDCSUQqlLG
WIlF8MVkS6f2POqFQyQ0JqKOTPHjGidOglLRoi0L6mWuhM9n1Gq3A7whC/5prE7QsF6GG1dl5yIh
xE/dn68saEQDKD05FOpmmcJQ4/Ao2ZrocJSSSD8AtRvx/X/2AAg/LHFGW0PQgxIZbgGL75UoOFq9
KNKitVVu0zQ2gF6Mg/LUhmZNdtoz+0kT8q79qS1PQRlllaCXbV3E1Wzz6gQ36eXa3eQcE9k2bQT4
KawWiHNZ4U3tXJLjgVyWL2rvylQPNTUX7SAO6COJhsTq61ciuAKhOzP4rjSdxI7fJCbKOLmQNqp6
PUamfXfHdqtIPzLD54NY0gnrxQIWUls7J7Kg7vEGY3eazZN/gMfO7FQOnSCDV37NnWT6f5uiNegN
o0JC3FuJcqwrWxpDMR5+5VQ2HtE3vpPf+7pwBfPUtz6WyHteUKEbnY+G7kHL/knLz8oJ4C0G85Wf
ja33gbhMV9V2QsIugQNC93QwIh9d1ihelRPDx8aSNYBiWhwiJJxX+nD6ZDs+WU07MW4JOfbNoX4E
O0j5XWCryKShi6b78v7GsAPbexmxyIA+EL6yr04z49tATtNUz7r6JY9re68TCQNhLs1Ck61ffz1D
1yWrIARHudlxQncnlxTGUxnLXqQpaHrQOmrhLReKzAEE4OaAWKYBvZu8ZIeNT9+eA1/lDqA6+IEK
BLwnjieXSt6F25b6paBinWnwKHNTQbUozj5wZlGk1hUwmYy61gaiQ8jL/Ifnbd3HVC+XRBx0uv/s
hlCMnEJjP5BawTHkfyLwpLUw8m/UkuWIK0uGhjxl8gwCV/EEMrBHJqOtjFTpgP/55oXlNsAs5rae
+CrOUrPItLa6uSCmReyxTVwq2TG29WxcIzPcmgDCa060uCZig5Ez698Irlb7VqSg/wpBWi37kNk9
zcelXyNdet0HEkj9BlFnIeJ8VqprsVKaYCq0fsdQ5IJTy9L/3CdxUehK6j4/tUE3KsYaCklEEwTd
kVwnx+xyaUIG7ks8Gzw62Z9vC3gaR6E724n+6QAU8+w8ZCxREm3Lo7HnlVxKMJSktQ0Dpx4GuTGL
JsboPkXY85+MAdZEI75SloKQmIMOBe0EgtJaubTyCvzaHaqqmmKmMz3HjkLzJXnh3THW+1O1w1LG
6cgvzldOmHoUbT45IDLqxFFz2Y58/fl/VEIp6NktsSmG7voICMGQqvBa4G8QhR/fXwz1AZ6phhsW
V6SrobeEjeUMe1nK8lJd+tDNKSOTCgphVbnO500eAwRmlW5gIoPePNMAVPzPZ4ZZk+/66jgcMeTy
Mf+64W8XMa7dvnNB6StLFqXZKjYKxB2F0X6WaCkPv0raqf8uRUYin6a2alXVsoH2YnXQ/SE9ZGSM
hlGxLwS+NuzTKuXKyV5JxExXEWN1Qlv9LHq1RQTRZ5B5viqUdf6Wbm3rPJqig65h5KPsY6gWxReD
TF80DxuuLS3FNpI0y0CaK4u28Xi//oMzkfHKRbcJw9e1sEb159OYaXWw4Ii2ND2pqE+eAW4uA9V9
5oj8E0JDw9eGAeecjbyCTUoo418Co/5+Y+Ioe0fcG9HY/ubDsgisv9ZLEiGwz+7eYYh3rPiWL/Xl
EhqmlK9u3qXgKbR7T30hoYQ9if2pgHEpOMlj3i/zuUa5N4tbg7Q/VMbOyrF7e2ZHuuas+JMjFWxg
TlF317dhodAggOrEyn5yszVXAdjVQEfzmgh36vfnvsuE2tXHUbMX9ApgYNVK1tlafDC/UHfaNf/3
JjMKbf8wcvkH3sBZpqCt32DExBvnwiI7icussLV93wtH8tLqHulEYQ/KMenXwGUmkMdoFuO65w9/
pBFr9VPqkFoNOywlbEij0Gnwaln1dPc5tCZzRJhYAERSQDVmrM4fyC3NjIa+FONF/yjMoe3Py6p6
GYVC2hVCqOlS6nbsCZnyCNiUTyNYFaDf/PkhzolMKqSfodmcj5ZSfVN/xlyUjRAwEdkzLCnhDEsk
8MLN7zshT6TfEVd7Qw1XfvvTMkwgEOCDGadbDmwCQGPXRJqOAGYi527ewaJasRc+FPNx9uaEBje4
ql3LSKlI7qCQdw9m351/DTIMTxgRlPQT2MS4CgiXuOeFCz6v2ht/GQ1rXHIIXAACMMK0lvORxLGp
8xGmKl1md6e21jg3qaFEKaLEt2z4nMZYjjnM4GE21841+uqHXjr7kei7dL28KPuBCwnRknooP/oD
TVfZuH5suOjojw+RvMcwo88P7xQ2kALmUvb26LdCzEDtd1RrOd3j4b6OUi5PQJ8QpppcERdOIG0p
ZmUaTPe9ZgaNIeDyrlxnlvl3UKFKihTz73vpgrvd4ta2tcG+1j/n4QJt/TdnqmaGfr4RX6Xx0AKZ
3+7Y/WcIngcAUKLMSGSwSRCD9sFLb9fNR7P4zehm0eZaGFPtTShD3AvBSvKJhBSRnCWtH1UDyXI7
JGfx
`pragma protect end_protected

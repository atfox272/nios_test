// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
vT0SE90OfFCicIVyP5y6ZYhZ0pI2DZVIYLxOB2GiUZpkTyZ1BAiYj+QyY5rd9jt7XGgkBNMCzmbk
kgEXT8EhM1q8YMiyV+QjK/5v0RrFtYEh2ctziMo/2Lp+W5nc7gxKPfvc40/IB8VhqIPaeeLrLECS
Nb0JrsBh2vNF1oI82yBU7tlM59FpkUdNNQkbGehLEdXN2i/085vAzfzIa6LTQwvtGMW8OdOK2VJC
Xs8zDlWmCk0AWenfTVoY5JF6TSlUvTCIuoiLijekUmLt80FSJ3RSKaNMVVxXYBzimq2qHxMF2+Do
na0dWgQ1YXcd6ZP+9KZSaRwYxNR8+3JyAYaXwQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 3376)
CG2M4oBJRr31+LqtMRJMZ/pPgxBxbjpvdIZGuT+5Mm8kZ3fuaeEqnoGaTg4v+lyp1ywPnr7eruWt
rHHZO0X62WEBTev4sJ6XWmTmVnCz2hwQE+r8bI5l0fiNceTdLcutOb2+m5kp7iVEVwO/g0pLUvQK
IusKL+fjhQER9jLzyBzBNd+OL9q55MjJPefqQHdMOcKHVA+cF+mwE3Ci2Sf/s49kBvAlYXI9XAZN
5DCy8EjugFOvv3t30VzKbU+2kU45Ttl2NrI/grJ+3CMcb5j53JOXrTM1FzWZZNxKjeB4uYXr4xa3
8Ge/N7nnXmWzjtOMNNcWAaWTllxOrEb4rCVNF3YYoUKkgJw72DLdN057RSdDV2sycTMquU1LXCHY
Q9bEAPcf+1FR9k+JXiKZj2drBWn3zKtdZC7t+oO094FCUnsoLXlZSIbIiBMhTQI20KPY0sH6tkQI
rjMnmxPjZD5et9bnoAWxtHLwjYv9kMIxCqQSRv8PawxH66tWbGMkhvYmRLb3nFuSL8Wg590r1Vdj
ZDA9cIePw0Q5JWZXxBesB7E6tMusFp/nr+H5EaFBfwvMh73urmOOhDOHXqI1rhqmQ5TZb9+WZAUD
SrPiyYJe8j10XNk2/W3bXoOBSdsrMbXM5y0QA/Ciao32f2/rolsjN3YNyJw9WL8pES0F+Zd8H5VZ
cE/IOrp8OScD9Xrc51Cxql9RLJKV0JX2ZO4FqNyn2qIfB74bWaMWtfKeOEkDu9XfrwBwP53jMsmj
K2oFWgbC3FMRX3qZPePLecvbn93zQhsTyQejleXeBq+wf3SdOG9VJy3TnXuvb0A2DKPMwe2yv3BS
nBcPOY9qgAyr4ZGoVctryGiTTp+f4ZuHsJpL0tsfkhxE5IDB1IEV7cW+sd7CqwsPlWlUsnn2MPYs
jCqWAGXUltbFFGx5nQF868RU99ed6kirzq9XrXVfza2y8P4KWWHlJ9TNfmruWNx2mYARI7Lq9PcV
GqAHyg3Ygtuyi1MnAfcheKL+sLgZM7s2pL85h16XtG0vRM7q+6SzuddnCjQm7ydqC1wRbc+MrRJh
WVQZaxhe3mSmg10Nvgm9PCmNaQJr2yaI+evwE/e4u8CowF/wye/ehwYUhThJlY8NXPVeFUdhYoa9
vFwrmCiRrqZaSLRTkcz014UaZhHUv9gqV9ANCGomHMrNPiE4JGYxZyJ4E9BlfmcgeXm+8OHl55tr
UpGdiry70TwH3pcCKqeQ/6qG4WnxuwT2srHXXl+LHphSCk1BZxa7fspehoBXPP14Sg2w7HzkYzlb
CZLbdApJOamNWksWDlazR7QIfOrNsuggEc/slq5LfWVsg2TqP3cUQj0V4RdVyPdkHv5UN9sMH5tq
Uycmbi9mhFMF10mL7yPjpFvey1Dx9msKEW3mkFhmVXnytOSpnfbBSDDYdklkhx/GbtxUPKW3XcIM
BLL5QVQPlbplT6QfvjriPH1tl+CSZu5lF+Uq3UbuWDMf6isZ8vyYF/8FfwYAmZE/HeSV+v5zU6+Y
rLCg+2hDjDxZr92A95grll6ElEqrb/yYdw0eR2KxK3sv6saQGd5Ee1SpqbizUhkaf1taQrZzxB4T
czhdvTlilAdg1nl3Z4SUq2uZmqJQ2u9ibteTs/WytjxFAhV8RraOI3zCUu7ckM93kRJssvypSXbF
4h9mvPUqeZJt7qnSGdNsjFTC9EK4EdXf4k926vYb2vfFAP0zdQvUVD82JO4V02x+nq+c7ZghgDV/
rF3zwfWWBvutlxV5P/zBIOVaPM+CeWbDCMGnHRY7VGqJGJSWpq6LVcKUKY20stZlaS5X6FDekjVp
da2oIR3jFCe/zMti7IrQkh/hB0IL1qEHMT6vGrJifjkjRFW0hS9XR+nmveSp+kh5v+OudFUK4v/R
kspMbQ5x46R/9KpA+lXD4TRWI9J6KlD2YhFYYXX4oHZ8ogVxw/PAj/4jIxKXwTzU+Hg0NiENWSnL
L0qVv+FXOLHqtvZysjgmPqqFoO25oAsYhyKyz+mNpnL2FBQcMNNJnUmH7BWLRS41SpVrBTRzaSVp
kzGu/2IM5jn5EeKPYqT7avO/aKcnijpWQdINsT1RkHccFrEdz2oXioXnbqCheGjfLW0dzXAnGuCA
sEoFYcOHoy3N1c7LdfgH7857ITEdm+ngRHniTZGssMF+h88QFDVD9FXQIonI2FscIM3b15M0s5ya
YhBawCzFSagSgQ+FsdMzWJwoyh+ZVJIYztO4Fr25cKfUC30paEK/cGZll3vzorPY5kpcOEFnupSD
NsWuHNB2WalRX4mlgQpRgz+o3bwYCdaczyDCBhCoKpnD81YbWvO1XzL1sD0SyO0WBIwFFWK0AXhf
Gan92o6RfLRLCVtqS+SgkGcg6PftFc4Zcji5gK96smkE3gNT3VYXIPwRwq35WEfZbxqtdQ3zMkrB
jhI4BV/X49cZpT1pZ7aPImsm41/c3KUvmOfL9tOuvRN8m95SHqo4lg+iDKTWh5urY5Kn/+RFYacw
aTYlhohHsJ4fi8XT2HGk2Lb5f3QDlpFV+RjFal7XYsxZiJB2uyJtKZB+4ygONd+1sDKLo2W6SthA
YhGuVwjo7vJxu6awpOBVGRcbAXHkbrrFWzKwvJolQx1LaCTkxhMqDdLcO0QxgKap43jy3tFUFDWs
z6etj39GLu1ooJw/8nt69MLQYiL0cNZ3QSiVjndk+08M9Q2aqcQ1s4e02yWLzqw/5w5hi0LP+3ac
cLHHtMRH9EJINfhIhoGWFkLARzEpyGxoRPk8xRB3lmGGU2rVWJVfncmVBBIM7bu8PD+cRobHBZtk
uyw8DLHcSV71yPynH/qTEff7d2gMeBHqntUv3NXX9+9bOmfZ19tOUtwz8fIkAZFOoY/B4/OpP3yX
vB9Okmk0QANVerA/BVPrGPF715/XjnWspNfVzB7fLTjv3eabdZZAM+yfzaqEcO3k4+3o6o862Vyb
7d5QVkTRBuu1DqdyuHLXn3lcx4E+wgguVXyPy7agnvD0iKZaV/PF0BSCPqUlzHdIpMI1AluHXobK
HQfFx4RVwFjL4glC5gIzdpYo54FUhQxEwsS1EK2mWwt0hRCKHoUV9RN3+2lrRaiUXxKwvwo+WyxS
bBwlem9c1rtCoM9TLYhk1vkOXfnSjNqOeR4Af4YWF8Ia3o7N9rgEhSi3lQcBW+MltKymMuGjZyRI
tSWiZG6z5wk0/KICbawsoE7/AXYW09//03rZ2sVrpDvlI2u7BXCO+oV3rs0P5+4qmA/xAFCCepjU
1IWnBUtRsmoDrn52SQOSd/izZ3ZZx6gNnCTm7Z/MgadoR5RkMxBL35VRWV/G+xo18Hp9ZvQSDfQY
b3obuXKLUROyBaIR2ZHylCyw0o/b7BfjVlnU5O2Wk1AbVUSl5VwGeF1sgQY1EMEpyWOc8ljy7qn5
eMfVfKmZEMbzfp5W9kbLlwyunk4lhgGLj7D8TNEH+VfYUAWs66iShQb6wvVzhLI7uBdliEsdb2mh
xJL8VUNCk4OYKVFl2biNwkJ07pAjEUDZazRfBT/uPnFIob0FZNzXzwdll0f/VgnD2pTQ+yTV5E/w
fkn3ppbeBPsxgb7UG/d0i5Qrh5pbHLos9GAYTE0Tno043sIQm8yY02kecnTfFeWOfqFQFdKiYOTZ
BUWWnaqEctpGJe0nMTedtv2kaat8Z3N2gc/oXg6TidxFe65c660y/5q7MSwAr5k9liiUjUwanq4f
FWOZ2kPY08vodIRTD2nkpYIZxjymLxiGYYO7to5Sk7GGhlP1rhluZwK1l0uyH1mhV+v2C5lp+F+T
qZIUFfqwGip/ItrtzVEZ9gYUG/B61Zhyq6JCpH0Z8VHRZTBn4n/11oanjq/kQNsQjudj3z/RFUlC
CWEUnNrpiHTdd+pqjF+WK/EUMgZsj31tXQFN0rLOPfmG54W/DCY6EyxXQbunnlh99x4jB5QbtsK0
v8QenTbOA+AvpOhPcL1YjKi3hPAfH5+/JX2sn+sxoUxVxSdv2SbOhCgGrFASPsb2nyXkSSu30Czq
mCC/LQ5DJuZWvCYeemmVoZ//OUlieNubNNRZdjvoVJOVA/nHvmi7Cum+Cm3Z4wM04ajauxxA/i7V
TGDsR5doqbuM3B9fYVkGWhnUoeY2V+hHVZMxvSnhOooJ1bnM5dDm0m3+wpho7VjTjmE1vbzIb/mf
qUpgg6WpbUjgX4zlheBMN0diWhVETeVsbAXhayxOJsu7sOMqJZxrpfwp1fkEsYcqThsbTMiK5YI5
68ltcC4lufh5Xs9yl0X7oDLTU+ZelZ1bazFiDkFEYxssI8jnwJmkigJAVUIkGp+2HDYM2Z1clHFm
SG94ZAtMLyfMqxJ72no7HZIHYws0ezOLul6buWuctAe1us3WR9enAiA2ek/s8iwDeHBZiSAQMX7u
uJjthRC8fkxTqY8PvhuqGWEs2UcGJs36erRR09V1ucz2wCbznJahj6emG10Ex804vilSA/RzVZ0r
MYSGNwMjuNJBxfyLOA==
`pragma protect end_protected

// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
RCAQV0gaxYs1bkb6NOgTrvm2z+WP/qxQJ+S8HSUlZ25GHe1nCsaJ+olKCA3Qs9qPXGrEdr4nBYnS
xrgPn3ixxffhkKS+tGoMs+HX9g8Wf1YIsZhZPioAB7oOODc3vUh693uzOOUyMlc5M2VOs93vJeOg
w4RZd4NvTa7Umn06wY9bX7UR5hRv2jA2+BXGvJfjZjg7Fpy1uTDvAdXucxEDBSorf9ZwggbC/hzp
/LXBok07y3LFIfkx9W4ddWRzPzbUXz2zSh7roJCsV/GQXy8R+SZt6AJUTxBQ2tG1pystKQgLrcoM
HDndysMMGDqKwmvCJQh6jz4oo2yQ3Crrz0DNxA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 73040)
5cDYlSKJO8VByLRQTaWZBgQrPlhyDnhPbL1PlkhdxUe3779vfKsYmIq8a95WYz1hb/k+XoLKnWOx
Cae3nuLseqInn9hb4mzYaeBjZIhmNyRkPiAjVeUmjQkuffTBTZgW4zIz4z/K0QntthJxwPvA7Aww
3DEdARtipJn2S8InAb4YCdKiGtHAYfAADgtLmpTsBUtY0ajD5iMhE4SZkNM9J7+qaWQH1plWeMKB
Xo9xV7PkHga4fFd1NmcnYh2z5ltkiXouk5Pt+BKut7fwGoHteHt1A8EJVjaXTDJ2NW7mUdM4klrF
d51zGUVE87WduK/gaNKcmAFZUwdKDt+GF3RSOiRAZc41Qy5qxjA1i55cEVyesHzA13MXbuinX9jv
3l227nVdY7jkpTy2MREsTs1uKgaDHpBWaMGBSqA9fBAEM9Pl2kx1O2NBsU3/ZGWeCiZZcciOPQKL
AIJnfadCqzLdhGd+Q6VPC63Wt4yag8dmgiBPEMJmDyy+kr4BF/UfKBLWOCs81yBAAuObcv7GnhvU
f6JkowOVGXWuys9lGVtiHk4jR8QLC9oaSyIY2XjjeWu9UImVr67WeXKFmhwXgyliTPj9asmeOFEk
WA6spM2NQKpr7EqIaPmrgW8BtxPsJevxn64IrvXWh0mhxAsM1yUxuQn/he2FqIGFP4DtO+LTZjDQ
0m9Gx263ArZJcS8HhCYLiK7zlRpGDqhGQeoFC9Ofj4glTvQ6z4VZLPq6OuNOeHO4Zj6rs+96ohFO
CadVzy5CmwSFyH3g6kL7MUF6Z5UnUljdLfmZ0jhwHX/A+l82yDiJWttexaa47SKs/fx+lX3ihsBz
XD2eeJO74mgQVfpjtOiAZ4f2HIwOHUeNv05NGkKfJgmlgDAdtJ7z70dfpslClkmnEbxGop1A8q5G
kZ6icZXuOtzgS1XNQ5WLLipYVkuFQAi5bzzRfzsZK0K1Ec2PqqtpGnqiK6FtCvXwMc6eH1vJ47c+
Qm9xd2JvwEMaqGHrQkmwWh6M5m2EdS4fOtjt2WI2io3UCSCWURMBrrMJV16zkalpyvafXMRSnHsW
jbStgxh4NOTCdCkB4bOKUjpy4jW4SDg9sHfQT13VTQlFunbHGhEpHAMLqRR084vWfFXujx/s8aPm
d8RlDQUOVgsnt+x/DRXD5mP7uA1I7wDYtGBCTAG6cl0TkdcNDiCgEqCeF/fJ7lVVzooCN1s8JlD6
7FsaDoVz0/Gzi2OKItBLL1j0OxFROsNyY+VabgBoxiET0Vdx4LwhVuiw5msTjP6ifKpVl1ZGb5YA
VFjqsl19UPl01g2neNIjnl+sRv8exfZyXrVoyjIlD819MUd85C8cqUT6v82fjtLf3RYpzlB/texP
+jHpaDOLcjZDTXlaOJS8/5a16E0KNRG7mK2cmqKV1Abueulumg6YCaqJ9SDknZYFob0ye4dW8sTG
O+KZBJ7+0iiEzp8T/jFZOcRlPE3fjRny2ePM7EJSqC9VepHaYDI12zBA8XS9Q0xMpI4tnBaBCzEg
A67R3wZbDH9f/RtD3IJEY1XuUlhpmQa81ZepbSjCOyAcatESmqVqISJnfum6xvgS3rld9pqS2PkT
I9b6vwcGTY+1qtvN1WYFDeJJjzKbfbdN+PqY+/ni+1rvKefTRi9dcr9BPmlBsVmGUlGB/lU9TNfk
iIx1xCH8Th790arMScb7Pl8YWQw8SMTOip4reL95zQgC+0UH1aiLegO+06yP5szOCHhlPLucJJh3
DZE4ujt3wHfHHjUjmQkDEBAmS8pQDkUI/bHU7Dq9yMk/XHmNeRJa9tcCgew7hd7eH4MBV+v9co3P
VJjyKcsJ6XQ8dxl0uEgzjT6mv4kpAHp9++Aiky9jY4CN8fMSCBD5fYqztkCn9ds27R6iaDyEC4rF
AFiIFOHyjG+Zlg1KDhJakFxIPQak9JA8uiX9uUGQa6IHPbzrPBtqQjRMzGCMyB3Y4LxXVG433v/l
YsgNnyPbVs0WxPR2ign99/PZrgspj5QLSEDg+9jW2GTN3i5HhHx4NW50F0KtCZp8JpTBXJknqdM5
W8/D4M4brRQtbR8LwwCmwrUNaXarR4629UGcLrJLhgsvYJHwoYW9o0qNVApyELU/vNon34A5pG1Z
woTUM0pdzlqGcgUf2U9XAiN431VGOBvItXorrXsijGxEigNPbeqbhs0XS75MXzy7yLPdRQVLLxDX
ykUWnKzDzUCtZNdTzrqoSCI8ciE6utmwD1kEHASzY25YHMAoNF8ocxcTqrjyPa6mMUAv2cXS7Cma
YSqzT9r1HAu3UYsOzvF3ZB+XiV4h9Os2wCbj7ruYBYpE2A2e0VlQhvy9nkRBIT9nCfdmLBBfZEY3
uG2Uk6kvVc0R4wb25p/l3Zuq1IAckeEtleFobvxSUsQ3nwfZVGFCR0zc47lGbjysfMXIhscP/6h3
AzTmOcZX9goG5KdGuyCwA5uvPyyHKs8tpayjDXDriyAgcWPezui3BswllGgqVvNFO+MaG4SCfMQ3
BWxvWoLvqCC00x6su+WtM593CMvVrf6XnQew1FUgv9HsGj1AO+jJy2wnQTEMuvGxAvS7UZs5DRq4
oIdISYz/go84z/U904MfyLE00AWWWb55QwgSNugqfGWv9SvFDPq61wiUzvD9mDn5WjXIxSGMsvlN
NpWRsR8EIZEN1juiNf48A6dXNdDEBDBl0K5JZ+13r5sIl+95HNCjb6BXD/e/ifbLIFgyz3/alMUT
g40lyvL9iCCleP+dIu0AG2Q6zdzSThKmMylhs5ORm2+gX02xKdbRrQnRmDctvzHbfTp/v8WEv8pO
HqePUTIXMGAHrAm0F47qRxMRKe7wySrjf8wTtbrhP+CZYZO2lFTwZUOkuIcQ0mfy3/jzHgkw2Mp0
hX0HPr/KorvUkzUEreUjYUOwF/mdYg2u+/nA7ve8Jg0a12E+SCbvZqf6dMjrqoyFl7CKRR8XDIEq
cQ/jXfDEntV/0FCyLItlT65F5+AwlDA5VC0WpwG6NVJ+Km4vvuGlrsZB0vE81dUnBEpj74EPa7lg
j9cE1LG2oBMURc5jI+WEZHZojc6nr+od1xnbcr7dmVWxEzVHFSlIQYq68ln7BOHU/kYthIz2TSsy
4IkClSr7S2+LLvCWJiPv4CoZsI1pH0hUzmfXzdahKymjLt+yWq8l4OKxFLsl8nYznEz9TN5+RqnY
CQIQx/20W59uyvtscgm/XnI4mzfePENhen81bJqzeoT74eFg+xHgv6HYRjwEQQwhSfIETMD8nM9+
p3zeS9IZR/7JGiQYoe3/0cO1g1Df8hi7XLiEeLQN62mnFmJhoPTCkMde+n7K5f8qAXD9keyk+PqZ
SNwpsRrTUmut276QGL5v1FzTKbyrjQ9uLK26c+zwHBJTic3/KgUOSHsmECuBJ6VucujKslSgfH2J
p/5EUsgO6V86iyJsbfmJkBBLvjqGaYKmiKFXfQG1pJawhiqCz9GCzeuGd8mces3qzlkybEvdxzp1
0QkNZUaKh5BK0azxXny1WjKKGAnYgHxxDS2FIf6KAVY01A1rWR015WDLGRYKjWshtjS1FPH523EF
8QVohSKsfqoZIQ+DxJbKcwDwnVaMkIKD2QOK6BL1Pek/99u04fxlHMWmi+KV5KsqXpeJmmjCWnIQ
roVVyiHNnqd/5F+tusyd1mHYtKQ7IC6Az0Guz3J+/pCYLHAR5ZgZag4CA1Q0izJE249k2NcMDsQn
PbmaKZtyIckN1DdK7JXkXCbufaeBnGcMCUme0cU6sGp9+ChgqyGu5VdPK2qzoFSp4VJhqeggCqfn
Z3cwkwANbGVsPUzBgkolpYYn358BV9tW17dKvCpNJLYimerHvDMqiBuUljq5KmrPUVcV6T62fhMr
Zm5ozYxmPVz4xm+24mw5nc+K/NEWiEhp4dM7plCB5EbComrQlueQnAr9HpLbvcygQxisHp/zA0F5
0Knu7Oh5g8qltRSDsOdt/+Rj9Gx2649b6hPpOQthlsratIn801fopyIg6Cd6kgyanpVLVFtwem+W
wKdxBNL7BIjAMugiWO6D9SfNNe6qaYoBknzE2FqnoDKdEukcxQp0pSn27s5l3gJOqbvM0gleREgL
QgKwVWwR3v3DzWFY/5kKoVF5cCLMew7jWvzL4Dr2nbGgyH8nxtTCd8ho9KZ2dXNyL0p7ME2uH+dn
FYZpFCqsMEgoIVxwI2XVj8+1ss4oQYO6JwuoW1CR56r1ZVKfDSaWaysCVdy/Ok8IFmqyOj9W2d8b
01iVhIGlhWd28kXv6ghW10AMu28j4fPyLX8L1kf4qTZKT+Jwmp8fMqQQ+KPcam4oPmQjIkal9X1l
ERA1/ApgygfCUI+wxcrecMib1IgpRcc/z3PartwyDyBhjCxHTUMV8Q2and+fdGwv/PGplkWVjYsM
UM68YB0NdS7QtiWOk+TmPKcEt6KRIBx2G06txI2MOq6HuAHs5DliUfpkaJr+Hsuk6c8InHGy27qQ
KL+/TbCQlm2bH9tnlMX6A+L2BWRQr4koIiQBUxHOJo8Q144JJz2IqhWBAVvCEI1DB+rScysWkI2O
k+0nkdKmUhyaK6M1TBNZh+eb/RV+Bol/2ge3LxEiS8wtHAieO4fEGMeR8tpkntr8/ZZk+tN1dMDX
h2OpK+1PWji5ANQDUs+Li1lG84G2KF8Sl5kwNRwouSNxDKOBZR47dLmKvxIWWCiyqOQGHJpaKp5q
24vaVFaMrK20/QiuPzVNohW069B7JFgd5n1P3jWDD0Fpu/iggB36PDTeiqzoP7tbsW7NEwlKY8FO
qeffDV6umuyQoWd+j9Ca6+M3Es6frC9p9wSwEMRdKmKyB0PX/g4RKgCwvGNwwug7y80LlNb7w0hW
Iu1yEUBMSCQQbGwcRvZg94tJsblApKEp+mpFxDHT07gDcU+pliIYMomG1yL3kFtVfPRatUHjurNf
d1Dpl4LV9L2wNebZfqaX2zaUpRQ9BCccvJoFo+a+YXQWuy1FwGGxG6le/cvf4TuUgvf05XZ0CH+H
h5mPY0GcQ1LM//TAips4bJ64GOnIbfygvnOiJxMn508dMwIN0cu3UWCQidWVxHpHsrWcqo23wqPt
qk9RUWfa1BIABNykxlWNELXdqzbqO+ljGsTJHPoTdNDJLNzkjaGWc5KcAOCorRHX03ZNWNlxIVdG
XDccoXzGRx+fQkdeOCvkV+fRW0Zv6A0urnrMvkn75tnOd0ldOC+PpUbqPw35dRo6mLTBvNdSSbJT
wCXAFVbrp3J8fxo0hOnUosRQaKzzmnBalLDkq5TCRL+ane6y3UEvgLARRziA3SovjAup0h5XdGMy
otKDAyf65F0pvw73UTqGDqdkjPPLOX+IoBV44DGSNQd3b6LGBzl7Z8SVFEnGdzyrUzazTpFwWXI+
H1nHfqm+eRCzmBkngk+7l0SJk1x6V/OZZtvgOKauixFV4/8f/BHWXbX+p3FqxZ8MZs6TOOXr2GGz
+jbI8fx3CgRbhbsAfCgXaELGYLa4UcOSeSEr9LifDDFdL3H5XU6NsQY3AdWgx9mhuf2/Ltwz9kAx
BUWKqU7YGJhj7i5YrNMGJDp1NGxD3eF2cdoEAcllG96ICLvv850d77F8FhhWTGaej3uHooBFcylA
z1FcHMOUY36x24xVKlY8GwvsvPhAlPwOAlOy7EjKN5WYGBwwKX70uSXb8nHsd5wZwUBWFj9m8oH/
9RWxq2ALyOrsdzfnkyIS/O03rV4u2jxd1jnvaPeIvCGO7Ow8cckRQiyvtvH8jHGYb0Cbw9rmyXbP
HVAx6n2Tr67g4C8ap0b/33PP020G1p2pxBNGIniV7TLqs5Jgh8KjmN+UmxoQCCXUSc3jmfJb3rya
Z8/w7F15hedgqosKuzn3XEA368MLN1+Agg1q4nDsaqB7En/EdURmuXznj30iReAVzS/7OZoIeAAH
dQwTjEgKUdEKObCRjxL/WFzSe7TwRhXTMYSsusYdyBm1ID8Ss8ePZp9yYYazudZlQ413vTmbdRD5
LJw4vN6+qi0pAitr8Vz+iZM2xp45Zd8Q7J5KLI1H1TzZXIsfamkbPeREMyknCSTP10kxL4ctCivt
XtRm6bVlfRxhofbSsDGbjU0ONuqwdIEqp7FyNddOBSJDv8PWieHal6ZKYNEC7gg2JpI2zyRs6pBr
M1qer1PKibADpyCsiVLoq4wuQ42I/xtXkvbSfksa3ciHaANq0PMPw2pME/VI+dTPlAZpBlhOpexT
FWuzCZp4mwW8waCQcoHQikLXu5lWpr249lcVdRd4+RXi/BSjK/cUryXqRHdXcWlPdvbn+n5oKg8I
O1ZMDoxDl5rIZY+SgfGnr7F5XPNG62DXHzUYLMuDsMUoM9EmtzgzChPl2LpadViWmMT3xU85taeE
I/i3yXvlSm1yeB9GlMcMwZhpixdirtACzwPfqHyjrtmplRHupR3PQB4KUropLURP10gdHczx9dLZ
RowO+pt+jYlHrcqc11Tfzrp+jCStyrhudCX0B95jl1mzibQigsYM5tcxaPA+CQ+Dc9/M+1Vfqgim
EZzm1nsxw7HxRglbMme/BcgT1+pppIZznAnkxt0ltnAeyVp2+yruPZLJyy6OVYM3CYIZ4wJ1ZVvs
xsWd6rwyEeIHqt6snekymxBpYHTxKak5VESEKGFtvU4bwDoOl2GYxkLroV1bnmAMkF0AgsvWKmLc
bMmBE+AINaXq4jMcO0dcS4CM2vPHp7IkqNUC/d2S1MEXxfFPCM/BidyKlRKCb3eKpmFqVR9BTcFH
7l0Ol8cXL14lZDwE+CiGaWJxtn7p81S9CCUqqOPTl8lu7y1In7NfAATu5z7bPznUQObGeSX4+wO3
yc0XbWVyfKMwkuLttENe6YXEHerYUUBb7zfqgVXjrq5wuOetv+B617LQKOBrsorvytu/ubz5NR+e
sps4EvDVHaEafQf1PByGhhRByvUUBHf1lQksmzFxFeQ9T+TVshAXp2OzyNvAWqcIdusSpBBCFTo7
S6XmHk3ChRuNaz/HY+dZ09MTZiIa8txWsConQb0iTJh64cUA6UXueNX2rVShMusPGALMaHJb4z7g
8WIH9lBCjKwicPyQuhWXvxlBb+lvFYA4GNpyHu7P4+MOVLQsVCwSbDjnOJfVRukU9nEGjCF0M6Qd
brGvqvF90V1pdw5OpcHO6UcQy59IPJumTYCpWnbYZTDs9s8k9VGkmZ0VU4qG0QScHZZU+keyX+Lq
oRPckOFuhVue2lRZVmFkEDan1ylLfX6g2kcQq6YvLbznQxyMNTFKfdBBraTW5yIq85mc2eTzxk22
tryv6vBfTqo8ip1HFmRkNKHvrKMjT0KALGij2t0IJ2wEUNDPGf3W7fgkTqSEopxoE19Vi5IguwDb
xZ1VeUmwW647NJ0wDnFvgYpgrJK9wLebu0uFJRfSAQ5uCmv1FVjKVr2urjfCz3d8zNEgPJAYYrIO
tThREtRRVOFPLzZr0bzALwaJFBSaGIQTAqaw9pIzsLWMSjsU0lzTmpsV9r9Oq2lxp4Jz9ozc8v+K
ao+i8h6EMNqX9+G3nwGuOlznz6aaV3Fpdi9WqewMEfCBrooeavaooYWRdwhP6xzxukJqe1Xb2rI0
guAObRZL8WjJmxNJqDqI2AKDRWTRmpwAl1cn50y+zLdcxDuTzp910TFcRSNtFPG9W/hksUDmFy7Q
K8waTfKEvgGDH6mfC+n6K54s3suWSJ54neeWttjr1lozNbVONNRTdX4uIh9Fq8qyCpuCld5vgrho
H/0dMdZQS7zYmqEX5DSui/uwA4Lx0mefpOuZx2RFPCSc/VMmnevjUbBNjy04Ovu9TCjZsSQ5BQsj
f4Pk0cz3XbvlnD8xRYtG2rSpksEgJfJnN+yE/ILYsEc11Wj/8JBBKPGh6Gc71ngD/ZLvgl20f2rQ
qnHm5uP/b1bkv+P8alJlPz4ESvzvRZZMX3/SelS5dusG3hN+TXY3BhN9O3Fnzx/7pPHHTIE4P4fk
/bd5jaAZ95PEjf7jkDn64db4+f/EgsbDp5z7D05eOKAutEH8QZGadQA77PWg+R5RiwgsZRcb8sKz
KUcmZFY3T3znONds+W2mNlK2F6gpA8+mwLDuXb/Ik4bfUgx73APIqxKCagju7qLfA3w3cT0UCgLt
MjC+QFhh0sw7dF/TSkYuTbND4Sec+RTR/b4fa73/NXTDlE20MLWnL5PpU3v8mbSIuzudbzU6E1SN
lMAiQaQojEhzw1oh13apooqM9W/sZRvOLFvJyGPt826YIMadOVsh1xcQvfJuWo/m4WLM5GXkaf99
xzt33fkAIafPLIGp0OivbTItjqiOfH0ms2KCi7iEwARnLXdY2Qsrqm3w652bEzmv7UL8s0AKibin
DC4aGmRygnJHf1U4mc1sHmAFbzMmHK/9egFHWcraDxNWu8KEVljvQM89KLwmtex27OkLQUTKIRny
l4ZM+4oj5ZE0l1ILTydDarboAigT1PhP/K5Z/Np1Iyhc++B5IjHEuIsO02VGr0fKKL7hc2z50Grw
jrG4TSzz3n8V48b8d87V9nj+WO0hICQ0oD3vXbfx6GgZK0CG3Cc+sbeB22bXebHg8mQhqPferfbW
Hh7yl+KrMpW2RZHJpcFrKkrK3tGiX/Z0f+8k4o4vF43t5MbHzb9u4V3nKipipYHgjxE/3iY4LKc5
Z1Cz789KNAlWvBqYUb9xA5p7I8+c2mKR+N8/OOS+SGETAcgwrLU9POopd/0vm1LI5wN3nYk0rxV2
6KBvo8utGy/qzT3edMfB5UEKceqIOEU4Oo8ryDcXUOvRUjBJDKypUXPkUPFwmXfeUDRt381V+wva
8I6Xh2r26d8Med78BL+10D/q/pk4TnVmjmqGI7OfbvOtzmrsv5vWqKMSyoughiUC+X5RfOEx00nV
iibn37LEX7tTX6hAgEQ1vc8MEuny9gb0KpOkCFpUN7fGWtaPSFYEzOJacJfNd2kJ09RjNypkdmeX
i8gHUxT6PlaY/X18CBoL8POgogRpi2Kzhu2ytaIRamCsqy4TnKuxCWaVVYioAOlJLy4tHn5LoZ6l
s+u9UJUU9dxe4rBVQLXkkOq4d3HcPzwFRGmjoMQr5Co4MCYITUtzIEH+mwBmHKepY8rc3z/dtpEo
t8jioHVTPjDOOIcfJJvV4TNTIF7RJm044z8z/J96gZD9YoYaSnUgh1+nr84o0XKjqNIFFvJaHyHq
TQhivnRuGUgFNN9FYb1nx5tF7qHn7u2b6saI+6I84WVOGdFksun+R9tOWybA7HHIqH9UU3mF1b6E
w0l2AAeltuNHHoYA6m/0+5aIH0vA16KynTRvsWv2uGN87wyazDa8HEHlHfV9lQlp7PWJcAVs1Oya
b1TWxIpp9RtMAGxa7vH5J7cKGeAPDZMmoWTg7A7KQyCcZ+7q4N2pv5JexKg/LSjxsAsmuqwsrDhZ
dZyxYGMjwzkJl52083oE50qrFYg1s/gTtIQtcDjakVRwEhssFu7T6fAIaDYFZ+Bl88Co5xQf1rEN
sBUjHhIPzWFRljru1THcbHNGAZp7K0j61snoG65h+JOJ1HDqfkCA8W5nHXxY9gtJhia9C+Q5niUC
wH48bdxISjvsGy27OsrzKo2dKoyoJn/LjxSrBqjuVN/1mJwGvNOMPEj+AU/6UK9IbxTOufsnF39k
LA13kwOG65rSolvsnqxhuXu3PVgVXgRyiRyogMD7vNOVN6lHYzFXFPLrSVR13p27snUkSBjNcJhR
W73VSUJ6agE4lnwDkVgXqJeaTu2eSfGIorFGm24hYYJkFiUHj9D0dZc2Lrjm6WguQ7z8Iez6Zx+A
WxstmxzM0YaxcCZeyT1BClgxPjBfgwe40HybRFydSWCyyEtVrW8Enb1Jl1HgiR/V5xxcDfSN/eAo
m7uXJEcM0kNKHfRXVnAjCq59qNwtT0kWWkVqYpf+mjn/JR5J+nKzGq/Uly8jbFcHm1m5/5cGoN4Z
RQohc2qpLIwybGA2gbQgAoCsuvWs00pd1mLAW9Sz/MQ0nITJn9i4qBfctHRWIfy4xatU+gmPimI3
EQi2hCka1cJSjS9IWVxuDHFbzOL+IVu7EeH+u3c2bg2ipp8NISvA6Ht2fJIlXsnGdOH1fKnFfpEk
V7HoOIna3/h/pp3XB6g2lQhD1qywRoIi3Nl7qSDABsCfib5LOKRDpz9X8wDO4vNVa1ZIlc8ZBcca
v7lN4rGuIskIrja1BB+7xi1fThHREF8NQAIS8Qig5oSoxhjIGmxXKQaMn4AuYN3fm5bd9ytQVYlY
RB3tO5JlDXHl3ACMwfIfYE8XCJL8JzgNSmR31Br6O1bmFWOWeiVIIZZzUk3KvaXkenvNNYNUqSlo
SVwFy9kGAXEsQ36LQV904rvdCWJBJ7NYkdbfYn7AmN7Njrp5yrmN7kSbecWgw/a1TOFa/RvVJZC/
zurpOTIo3cC1i+IB1tCWRlBv824ps/9NI7L+8CL3xOd7APLwgCwTYIja/FHTLPt1ZPr5EiD6qN3L
zcCbBbMvY5Kzh3Ij4qSVyfYTnrVPo4g87Bx2QAQ7VEfYM1PN/FSJuRvLbSo4fR6rTdxiNUtQa+Gn
PC5yArgYUSokY1+1yThtyhjutt5VmMAbNEGjtcqnvFAowHu9fMEEJppyfccdjy1tiDjHt34dOuIZ
YpesWszwN/KgZ4RQjTyAGbcvwQoNjlYwbt20h+eMFO5jqjAXLve81eLS1OXqE8T88PjkBBddYoCY
PTf5qkfY355o7H5YE4FVxzFUBqZpaP0OGXUu9JJAFsRrEIBkqp/AHDnK6gXhS9P/ArSDmj/CMmLQ
UBofG5/ZlZ00XiIjj7C5IFMgiwgADut8VwqlRTzMrZGWXjEd3BHbXAOREEYL7PqH/qWTNJ00rTiz
s4WA1gEysBzQaJ45c/OeIj9WLtdKiYC/X1JjJSbgrCx8PSI8WDGlcZk/hFIzJqsFiOOl864pMfoU
OmKQ5vdcVQgrXrTZKDfTgZN0GVEwAvBz0jZefK2NNVEjH4sqA7nWTjFlMJL+Zp3gDanxTLQyBOHr
3B6xdqemJPdOJILHv/jrwlfKjssPxuywUY9jKqzPcnthEyd29IDClqvXi0C3TfVzbMt7D9jQrVq0
7HkkrXR5x4D3mUJILXpL0oUPZwVqAS5/Uq9UqZCyGwZYFZtnfZ7UdFXOZ8sBpdccphDysi0VhGy/
RAkp4FycnhnMzX1j4FtSmgeOWS4k8I6Tdza9HLircReohs7LDn+kP2SGEyLLjiA/7UVlzjPVY0Az
lzV29xwxYD/76Xb5zVv1qE447qRTnVd3I6Iqwo+PihNG4IEyTcblw9IgQtW2008iOXxvQxKIblam
fkgb48Dja0fmRXV9L/lJwW7k/KnCEXvchmcmV2AsvZdFoVbaZDrn1fia+tXspJkR2ibTxy56+8px
l875v7+yarXIktA5tkXs+zx3orqC4VFjQGkHVTLeUEP84hr5Vtq5dnyvazFvqBMtNOm1rptyySLw
nQ1rwOoqvA0uqJ8uLP3n0gZMqiAyEwenX3ByTbK4S97+j6/vvPST0iD/mma7Q6H/elzBOk28M4uB
EhuHIv7Vz7bLLCHGx9GzuC5XDeAGP8PgYUdqngKcKkZXJaSSfueV/v9NghSqoYchb7MI6QTno+Bb
VbnAtgqgUWTjPjyL7d5NmLPCUYVZqvf+Rj+AHXNBqBH+88bq7T6ZfEQXykDtYLVoaCN98bGByaLP
b/NIDTcKizmsjTKeSBdn9PRv7xD2T/q3u8h32zs1WvFetZZ0gpo/dCocrgJWzjAeZcDeT7rJ9T1O
5up3VKuqz/5GkF+NygdqFqSfuYeGjn5OvRLfxfoW9rp9K2Ekhn6oCpUliM6ikW2+tYU/24BQ2dUT
duBURCvBoTDQnm3pHq6Mv3MiUTmwd9h65XhGHwn52tXoWtcfmai/J/ZUuAKQDvXIFjk6IF0yigIu
305EDha3nZyhYa3sKzDmA1HLSy39twuIlpyfBJ2ypHT6y+3+M3YQ8IOPWgeVRLkqfJSEfQvH1ZCT
WZboHhS0AShkxKp5/QTkPw55hChf2K+mMUG6UfdP487kED4plFMgpPeBanSFuv4Mu79oO8ekeNyM
fqSjWKGtyYIunxZ+mLQ2fmtwj2irp9AdRdfbJQ2YZ0vseA/xk3rMmhiJoDbs7jmDdWMyxXkDQ7RD
W3xYySqvaPzcszs8ly9T8Ro9jXsaE445XALkFKojvtOaJYufry3b6L3kdrSpz/JCuRrHYuAq9pob
CfFbmqlERTkNycrmeefTA3P4Q1cycGtuW57Cc8Nld11M4jM73ZpevsXCuFfjQhG0XTpGpygzAgZ4
tDzn1GmkJGzuabnYVGA6GhHSPuXd6a5g+cuIYMLUpJVjH0Qhq6Wz7avPPlxt9og9bpRgPuwT8CE2
iWgdI0PHR64+INbJwosSGliY/kOxI8+T++VyaLZe+iE6C7mMkG37EFYnRKQpqVWejWz+qh2lusP4
+8zhrjn4fxCXzBQGvP61FWCiuJ9yr5/7mR7+NOcOSceta83yevWULgXHZa0XqJuSIlVURoF2+QUV
WYcPhRzysSpx1sMl9xoUTnvM3+tweAh9TapyFy1objBFAkAO2J9qBc2luCN5sV3rYBBZClXu6j2z
EP29Q/+dojFFApqQcviMEadbqKQO3QEm+yrKIf3rGXbwQKI8+4faBfeB3+vzG0k0PBZ1bI8Txpug
d6GPfgapnoCjtp44z3neML1EJ6c8qkM+9Tv6t9YmZMALrtr8fsPpktmOq7q3XMb8TsvOA+Xm+2AN
vxhrENaMMupat3TLDZnxo2Tjuket5cirFRGtphgX2Aba6OZQMl6zLvJULY6kRZ6z4Qvtzi3hyUhi
5wn7Qbw8arP9JHUhLclJ0lpGC/zkrDVWopDBK9NntomuQ1AIzbnGkekf/XnbT5djqQyf4Fn60f0z
DXNwR5g647or8UHMxWtSNftcIeusJS/8ak+FqLnyNqOJsBunkQRMmOMARy7wO9n/sGnW55Uohfy1
qhXUKXkmGv6svoFRo2B+BC3OAa+5/H0w6ql4GGW+UZwVAT5qHKYr8vveoD1U48xgKJzJtzr3BCKh
q70F1aLJ/qP/85S+bKgQxdgVg+IVIHMSFBYsFNxE3uxyaOpoLAn9pv6pSirnFMeOnhjukvsafNah
3Sc5r3t7FxNB4husqD8Orsmuj/d4HJ3p5JMzu01saBaMlvc8IrIn9WQcmNiEcx7RfEcZ70CHbI09
g2HNGP6nS/WBtt8KNRi/fcf7JWRBc6GYOc+PjEX/y6dWlamG1y2176tmiva140SOv0haJ6Mjk99I
DpNQTyY+9RypiZREu55vjRnGdaVCt5fARlOwygUCAM3EGCHNuDxGmdVo/O9kJK7++7QMrpfDnhp2
gNVt5p3JsfSPq3G8cajZfNeb3pno/u6Lk14FuIm7iQpHXmFU1f4SXa2m6HaqBiWVj+Gn4amj1Z+z
zp1cCZ/JLhHPtpeZSvC8RrvXNTLV/VBaSoMi8YySK2noKY8sXRovBU04v6Gprdc36vnxPZ4AZ9Vp
uviZWOVP3VCNiVnDUmuHssrHzMFDsZjZupcvW/MX6AhzYlL1skyEcCdB6O3bd7PjLSYDX2kN+KEB
qpQdZGaS2Mi4pRaFIh2rHQXfa4aB9DReej3sq2Bpo8K6qaHnWSoRjE2wgfD7eesjVcrrpLKbXFU6
aXcxMAj6Iw/+OPreRW6qPqrFT7d/42Ceh1FbcSsHKHOenriRfamgF8yYaO9dBynyV2h1qWlChg0x
55wRVZqnnDRkS6tOmOlDwBKT9+lbjM2S71CPpgeo2nttNV0OsOvdE9JLse522nNbxtq9mIMrd39M
qOI0fOo7RrCJJeEssQ8N/agV+0GkMCuq8jbU4eA8rnzD/0FpRS8gtZemvD3cibsC45Mczn3XJV7L
hLH+kOyFsSRBE4pOMoLrLS/a7bsoxrzfa5lM7E8fdyk09+RYBwEi97wQPqP0gWPdX2n2hsr1+HKw
BqJc0hW0lvNABruQTOQXXnB/AAwi5/2rp8cNJM7XePNdFZKr9i8bEsI+CJkUtUV6bgsbjIMu74C2
Y2+ZlxhvLJp7TD4xlPRm+PKhF6/P/ziX0qzujV0T6SejsLwSjw/tSU2KBEb47fSUvb3YiyAtnhxt
yDhLzZaNdWevDmYVmuzbCRJSH1GuRo9nhqe7WQ10v8dDVb4VOCE4nUPHuq0FtPGDMJgYPIbUR3OK
SOtNR0mzDGSVsdaTzmUHfwXlp5WzdDMjaSIIsdq8yMwEOs7kSf5Njr/zXvL8AglmjojXmgeaXvUz
IIon5dWu5vF2Vozy/kpJ/US66K6ckQD7otauAglG8C+hA5yiyoDeqbdapVVN3vJSi7bshfOzkqGz
f8npwWnNyr2geFaR7Qb5laO6/cVegkS33Sc8cwUUU/hpnUl0wBtEj2CBBxY/FpEcdqFYOkwWXNPn
pYfVth6CfbWo8Gqei2eNAd2rPSmM+YEWoKEQFvPwwF+INiTG/xrUr7s1vZDG2r1RosDKgtVdXL3v
HZW6dRbybvCqDtJMU1ubojlKvQ+HlqNltXWc5AviLyqHaLdXmNgybcE7zjFROS8bR0GA3Kjqbsal
+BLgSDdjBr719zYC5xK9kOEI1Akod4E8/xENpHyiU/WTUvZ2zFdd5J6NzsfglFdzUYVSm8AiT/RA
og1aaoJ2aNrlgL821xExi4ZBvkZkEZ/FcnY2Hevz04f/rOP64CYmqCbGUg/F6ZhDP2xCsfj7SH1c
HMhCWrJSM3k7yrJhSbARXgiXdSdvN5+3nig0XnHTqlU1XhZMIYfFQ+UyR7VPZpMD2ZrCTfRj2YLh
Ou66x1zSspvamRS0C/xRodGbxS4oH9dh6B/chiiT6pt7Gh5Gs0rekGUSzp6UTo1NNcvvWOJqT4ia
44vWmuSUxdymgyrhM0Y8AbeIN/1dUjgdpaqyzuxzvwoV2zxznGg/E9rXYXJCPgVqmEuIdwm5YXVV
v4sv2HyiRqy7/MgfGarc+H6mSCUbHFvwf5hCwa4EmYEVsQPrK3mNiVg0yHKeFJ9OO1hKSXt2umuY
6ak5GLyx28W6lO1yBFlUp7bmOH8WnQ3hfv9a1ftHCwP+YdzH6eB3KyicSzZqbf0BGXZLdByDOPUf
h/r20VzawJ656xKZ7MP3RulKZsbORkNU44Yf5Xc7Iga+gWP4PgH2bgwyd/0MNKYu+ZCNn4Rzfx2J
TucVt3eWNSy9Se6PpGYrOjjl1X6uKs9A0/lnvpGoU71mLuQ+TiRNb4M3nWQsSTcZZ5ucDS2cBIlh
eg/WchJmRzp89GxXxdvFeicZKjlxfFXvBCsCJTNLpFkP87ztfJve0zY/RgnXQGSKxytfZV5oZ2Bz
muFVfnJYPIP8zH0jpV2kLJkY3CHKKxjeWh7WUmy+5CklhUAJav811UIkQS90EJw1+9ZFDnU5+tfm
CBIGlK7I6rs+KWj3Ow3TYQ5HpR6HntusaFnxUsS0hBiAUpdadXwKFle12BQykJA5E941V120S2Td
V2C8YbZVWdZ3sza5l00FvU1xKro4blyEiO4XRpBdW9ZkODfqAyk6irbN7X+oeW8wJWpRotNcN3vZ
lsyhZBABESm7v7RKnxZwL3PxCJ8AndS3EXn1rBTcUz69ap1JcFezKQSpOCBi+uSQwlNdpeWOkqY1
mbwg8iB9edxikdbBEYnJ9GkIzJ4BXaxh0PNw+Xs3/s+77eyGDagDU/ZAjudEkIumtynL2DMabME/
Ppnnb9G9X1nJJX7DzZv1lOQAhRM/np8o3tboG+AP/w2vFvy/A0eydydyaTvJi3TpBV/qst4FkYDb
ayQGRAWRZ93MXxH3Dt7TDnC4rVmkA84+jrxs2wtAqy6hmO48ycYEenDcY0ewTRlZax2PHRkBuWPp
ilKWvs6xHmN8rq+7oMNN4huVoNW7c63fbEV0XBzHslez6lLfQPEXg6CcuKqWwTRrehHTozT5a1ci
PGChPkt9EcJKUzQuKMyJeUFo9XyniQShGmH6KNHEGae8zo5isA+1nVF56r2Uu4txbCTLwoyvlFOL
ArWROEA6k5XqdINkvBPOi1sIQist/EcU2g2M3Rc0f4xexs+D2P5bt7l3EJlo0rWxtRmaDColW+bj
iFKVrf+BW+HIE+AUmyOF52gEoDOwT9F8RxtELHNPIGCCCsRTLw6H0mhbpnhO7pVymCunby14rGBq
Tf/TrQvzfJnZq0x2zj314Oht+87A2zAZR0bqfdmLjqtYF4kNKDvkLQEYuCwlqaCPdovsphE9yUrZ
SjSI+XuUY7D3J+c5nDWNsOFp3H797+JYNwD4QNsQwOmZB3eaFYPhNRRQSbwV9/sY+jkOy09zxBGU
+7VsK+8g1tRdkAqz6y3LtamfScIuQQpSLa8aARzn4lGnv1AG1QTg+I3fae5amS5NoKC+eesJRHXG
H++NhNuEH0ngXPk19IgCy8ytG5HfU7ytIKFffStcTWPJ346XpoXRN7fQ8WWz6S1+u66JqCQJ+rAU
B70BTgPb3U/+tEP3MMvLYbXW1+rcK4TyfUYct+dWxCpUv1spMKaiXsDJBI6uKyM3CxmTbhjOomXu
1ugPPvkBsFfPxldH379QT4xGgg2RyQpomUfnOwVIvSMxX4wQqmrvVE3rHnTMeffuGtE5cwiPm7hF
huS97GGfctJvCRXLuaMuQvWA2udBVdbXTurVgIuN49rLD8L9QSRVAk0XjN23b2YJpp/wTKI7R7Zs
PnsPva7FySzFVM/uBVZOSt36Ud6aR/0Y3Fce07K6vy3TN11+WCJSOKiQQg3z2e6m3uUCO8WjeSau
Nl6pOPl+E32ydHAXxfu1EzlONyn5gXQCPZKYch4tQHoJNI9/kDbqKIRFtmQSHuvrN4P5hu+6DGEu
x5EUwmPZlC5GkBK/gPpeLRm7FFjVyrLDU74ZuE0VnA6fLTOZqj7Dtt8Ep02NTf4AxOF7VaF1TFL9
K7nz4bGGM6QEECXE42+P5R1ZZoQ/izd1fHkRYnhWR5CWxd2Kp1WxE41H6yNpPSFrzy1SKKSOYmfI
1kXU10pUTIJu2zBwWM3bZQJkJhv7OeBcdZ+RJTBlMs/fsXDGlGx4rXuaRByvIJo2TKOrpyIaQlrc
UUl8sHSWlWkrLrrZ8E6PApoto0Qaxnf2MPrVuQNt217U5Y1zIYTwnOjm3geMFQHOc2cbQMRtcyUn
WGT6msOBiJ1Qq3sNAMs1f8vWICQkfli8Jgtd5CYN4bKszKOdViXFPR+zCm7g1hojNX9URnpUeZ4i
N1f0H3gYBDF6XcW0vx3Z89Zk2745LbUzzxFnAAArlXfWqFLNzNeKajr9tKYgrbaHSHQDwnW14Vgc
p121V07i0/GeVQTQXj60PL5APwfMIYYzVFg+l0nj80wExwCKERp7Rq2TuOiUOSRwUwG5tPgXSGdn
ZZbx5JNjxv+YQ7QoqkUIsWXGEffqtaUwRgyGpz4B+gAYdazrgEXjJdfFoG/LX8B0s48KIGuXhJ01
i0/FEXPiRE8v+RTUQ71ATS+hFNqWk5hqVcQiYkwL+hPZgSosVRfV4wmFP/xEK/pX57v5RlqX57Uu
9EnW99tQVJR+v/mCpqP4VZTMC1RhucP+EUtIysiMrkoxByN78RHaPOzEDeCMYRJ/k7cVITgRt1qQ
TKbSvRZMT/pZZ6VL0FQrjHS6xWklA17f9ZugOwhKargwM87fqwYDAaP+PIvxGvCt32rOZIbzYFmx
bYv/rIH5gL8irRdbNgOuIqKLFSpj1eHahV6P8GwhS2c6MkyTHzvrrcKZrVMPFJq9ehovs5wCIuI2
B9cVvrG+53oF2hHflANKncBWFrQS5g4I7QHXBrvRXyBb/vY7EjpknzW/woZ2vacRszIaz0XUd421
j+D4Mc877Lrh5sCyO3zR+ju3yZ8epFLWDstxWr1A1FoAST7eFPDt0aH//UbIdJWGndf4MvujO2vz
BoaeG3D9OjjJJaCIx0V6Vx1tXezL8MPJAp3mlMrqllRVXwHCgj2MGUGbbzeUHPmHaHE20fqjjn/m
A/nRfyeGWpvHGO48hB+Fa4NJXwQ6u116FV7PfZs21KCp0FFe+QXo8L7zj7973kLZ0/el+KqVuSbU
TFZRZLUQEgbOQdt7vlJY27IDiYg7NhwmUId9f8l6SE0VICO2Jxcq3Hl1upbEaP4dTwmKZnlmltqO
lFPo/D7gWx+fZM4W/IfDS+pieDUlonWzYOF2OUlUe1oLJWhJT9O79s4sl5CqqVw3/3RYSJ/EA1Bf
tDRWtujKmsNh6QOJanJKXS77adEpQSC/h+upo1dzf8An9S5JTBqnxHANRSeKs7npMVjs8zQzdgFK
m6JLb0Jpxw5PgCnZZxB4q1mn4caexlZLcxsO6W4PGXZn2DuJP8iZYXNoiiKcZSFGU48lBqMuSPFM
gC+TfMjmbv7v6yWUfjPYw9F7qXxERzk23g0QIAJ+sljHw++vU44N7DLMBSHrBgDwJtrE+3iDwv61
ccpnelBtMwJhUWkYnJpORvWCV0TqMFE83N6WOIosg/eH0stlT/Fa8xsaCkKFIxQ+p7A4P+SpRoXK
GiuVbLMVBnzQa51BuEyo+G40Olmmy+DU4ooQnJWDFyXMRWpCsrDyyQB5KDIJ/9AhbxXl5FVlATrh
FaEu2vwEDlIqdnugYiCeqqLEN5P87i9u0zbfQK+7/2fFupOI8E8Id6HlQyClnqovSvO+AKjaBWmT
jCP+Mcg/uVAyoz+bBhEWPUwQGPL7Ro6ubRmXiLYaOb+wZueEaLtySmNpsY8DYAsLMYG9eh+7pKeL
UFwWgwRt7ASP5TTe0UGossXNljqJXe2RAvGqsah+ZBtKER7UvsTDjlwpChSxrwhCoCiKNvRpDvKt
FsaVt8Fs2GQLTQIv2NFVvARFutcnqZGrPtSxs4xoFbzLESm+jElsLRmTr0oUB3uZNm1bfT7OZ2ST
PO9B6saQMvyIzHu7ljBTzqlM75d3cN3D8Zs9txejxYc2xb/MVx79Gpu043e+hRu5E2NeWpKEO6VM
1csh7aq5Y5IMZbgwctwP4tt3EiPouSzN1ah+hjbCwD1bH7v+RNjpyFJZ9G4T0FwxtxLqH7qm746m
B4J1csJLGgcMvoleZIEi/ORQp9jk7IDCWkn60O1pqtjYDt3J4adcMqLkkgAHoCj0HDQkoioRhQ6R
CF5iswh4p68/e2Ekycsvo28OFpo29ljy9CctM96cX9Uxq/jS5+jUugPYm/v55QI3Ol1ok6DCdx3k
osnprCP2HwM0pgvku1821jOq657wKR/2vuaLcSXQXl5p5Ic0F2njlnADoys4GWho827TYo1flvs1
s6yPwnMcnDWFBiGkmDe9d8czT9FMINGOn/bG/kUaSY8QH30viAzKkw1EaTykSmR7K/SDUFzMywv4
ehQTzjv2uWh48igQl0TTeLaGSsSbeYc/QY4hijNUstXGXF5vrFqXMZd6mDzkM7PXzXjEu5IBDLWM
teN3x1DQf+QAXvy5a2Jj7VVB2KfQ8tuYDwdZXlHCBsxC05rZREKgjqUdUnVh2L4m/EX9YZkHYeTl
0oo4INNuK6aHbUxG1uDmpPWhNSdqCPMJh9Psq+FnzYFJdz9wV3s7wLPJE0CxiUwgpVapU91HAXND
mertibRVcPnzm3nzNg4Fc9Az9hNsgqnafeCQVsoDetYJ6GkzwoR6Pl7Bq7ZHSpdCvbxYrY0WFkIy
olQheZVFHFu9zjIujTHAJJ25ibI5Tj4Rj34nf1bG06Pn/NmixeN2zairPY88gdRFmp+Nmg+2UilK
rGxTxT0U2TJFFlCTOu1x6lVjXw63hM3KKoH/ZCJfwcUIPVRCO7g2hjJGKg/cuFTW6O1j3rvfyS49
V9aozyup08ZIKMMRfeu8agCu7nlK/lmWxLfCehfkZMt53jDrvxTQ42iCugNO90XnwADdk0HgdA+V
sIIZUT4li3IuY7HUZxiXqv4FiBdxpg5MYHvvwnI5QNbG3BhvAaBvu+AbZnPguci5ATyVzRMDsrC0
tMcoHmUVfSCKyturC1sUEHi/2elpc6aXDIq7qb671xmEd7t/IX4IQRMAOHBYxAVUo0EODOXMCIX+
aFlodNOQhN6Nsy7oEhjIaFGzLLo7Rj7oMIz+MGdqBi19TSAng+4axhjoDZs0LF0HSxggbqqZlK88
ULYdycMLaumv0gCSLtVL7y8wEtTg1aj1cAAOLHOM+EiGhydw1CV0cpCp49e+osi0NrXi6uaRWGAk
JY5vz+9YTa4R/i/KSIoTSn4zj6WUi7+j+Va816O0vaeOeJ/WE+plH4vYDKUm320HQ1wIQpLvZExH
pn19QDKrwgLULSW7GPjqTxGtMzSyt/cQGhMvfdGQ+wJg0bl+4xOCsckfC1lRtQwD+JKdDlaJgBZJ
jgkjedY981IaEDpxA20kmZhYBQfGc1aRkmafiTBNJB8jf7YIEOqlbKlTBc8rlqb/iZDfjZXOxftL
FCNX5zLeRnQ5MT3BOatD+WK/vTZLNLhuoyvO8g/KyJ1D0Xu/WmfwCvMcyDIG05TyzuMV6bKDQtuo
bpXIW6Hn0opw3sZ3Xs/Rf2C1WUeXFVC+6R1w2mKaghN/xeqFlKcbLc5PLDbhLwUdjSbJyy34Ih+y
TQoH4BsUB6lpgN6oxOW2KpqkYFmSdhzW00kBFpsBV50G1vCONIDuSOu6Dr6A1hmygzcMAXK8rsO5
IQaOIstbX9XXfH47ku3r1bzQ4n+JoMyR/FDKy0H1tmFVfeAxL8yTCKakGanr7KSLQ3HIpHjAElGP
3657ekOJYcp/Q0m7qVXNqh75TsUkui6SZQh0URDoX9R5feYjPl07FmWmDjMx3TEo7Bwle88YS/iL
TmoNvSoakHNYxMSamsHCH0a7WNYXQY4SqwymTLZFdjo2vJxzl9N4zJN01EtWxoKSLteG5NYSswjY
HwwcasCTt+Pa6OxwNn4ZdRDhlyPwCX4P7aYy7RnlDgENBDnjvIBoAd/iue+ncUzAcnMUyF7snUfu
N03a3kVlrJLIfG51qzTqruzD8qn0vd+szF7pyyjtytzf9IXAd8bgQlNVJZHxSZyu3U8HkuC6dgEC
5nvkcZvO/FCp+1zIdZw08uA/WaG/QXIxMY+9OFqSO6VqVgxrfCCXCNqCadG45vrIeJbWJWY2au3V
1HvTM+sWBN4RWalijQwO83217Z9Om95pjDeGqVzJ3DCEFzrUe8La7l1PBwOZl74LZXY8Cf28xa3B
wRmNCF38osy9MHQXYYbBIuSn95Mu13e4pPFv/wSOQc3bZQ+JmtFnI24KKWYj8RK+oU7mUeKpCQHf
Ucc+Km6j+S5osDSrPCdqTelOv9//5WgEOLTNE1fF+EGmbW7OMhxOFADJQNqSLyFss0g83PPehhUD
vjBBQXtgOr2DupTuWolf9xCRV+2e3ZTgk03SUp9K0/ZLRrpPG8lSOoQIUI5wH/GtgZNFOaR6aOzj
IZQ2ekGDlc+NKzUJ+lF0xK9EOlmmwLwcPh19xmlKw1Ws+8ij6GnLrr+Yu9Vafa+G28hRMjtmihUM
d4jwnsiqPrd/RueA420b6NR1M0VwXKIQDIxuTUR3lx2Mle54w5x07d6jIJbbEqzLy4Gqz7yskXZS
Hmm/4RqO0n4bspq/tpJv+gPgTdGQ61/fwfsGy0rIi/cesdWLxGn4Sl+/cf9Xeu/HfqFLuOWZ/xbJ
xElNXDgiVCTYEOteTcwd3ueu2Ot3CdvQTs5FFxl3UYYzODkJthh5e7iZxxL8BdXEypRKZk9K1A3o
g4A3amDMJ/MHHwL2sjSBu1Bor7OuwDOyC9w0KNROHMPaQKX189T7jFRkUhQ6zL8l+GNnuPh+zHv7
IHSPO9OwAePVUhxhxzTrAmhmlhLJncVO9VNaWt1xsAB/Oo+sIZChALf3b8njOcit1oZ6P+2AUmiB
MS5pVBmU9FRid4tWCjx1lw8Ssbgs/AMETuWjQpX8sTB8Ke50DZatuKOUZ3tbNM3DsntcCYtkE81q
HorY2jX1d2nkUjhTKbFfbFZTFSAaWciExUyQL3PlBPq2esofoUBOJ+Gm5/h5YHp3dvM2V2C+7Chv
gQWP7YLhj6FegfPy5HDt2hkfz4fovZDCruaoC9C/4fDxii6jmVD2E5qQtGSqziqWNfH9JBsCeAdl
F5l7S3o2Sf3db8dRymqEKl78PUR3wk6115HnKIOYr+QKyt+nMzJbkdkWluJVfN8y7oCZg0SFEGYB
/xancAYC72eF9Zn8wf5Du+7JoKEmUZxQoN/wC6tMURCd64uRzWBqxcGSPR5tYNnxFVjHFEwLBM/B
zrEA0f8dtxdWyAUrAaZjwpr0Vj09Joq44xgZ9eDwcN9eM74a4sVNTIOQu00zs4oI7hYJGiNPKdIx
v2P1nHAzpe+0nPyp0ioS8qboCHMjeTdQsAe/CpQ6S5AGVHlUerO4DVGJxiZoZ8VCzY78sytSM5s6
xkLesFP48Uy+uRVxyD3EQuvIoKeWkamiQj3AzjK+PQF2CGIwWzJyO49Dl077xxcAhO/jhv0YMTG0
o8qMJedJGxDO+VxmodqqlZkAn0+Mci0SFxjXFLKXMfo0VjQNtFsUv9WFCs87ROtdgEjLYAvcdNTQ
/opbzztzqNhWwfwftz0QIE6MRRlLw3QGNTRnu6xdkf6lzZeh42QNMdLQbGU4opF359YUas+kKnr9
n0k8rAOA3cizyGRVo0bfOtljXmif7Y5T00FAb5FVATFXHnIQOhg8QY1fbcI9VwGAqjMl56Wx9/gc
70k1YPd/M88A75OZ9eEJzVa2VALX/0TIeUYFh1BWTO5CDIRah+N5SUe9Kvdc+YNkP+paMRQK+2ZC
uXiXCglMadbClGpGJygN3EYyid9EjFpL8RuCdbC0rhekKOV+tLzbEnp7SfJh2KlIDXviN46XXXcm
U1wfkWXDEI8ZtwALwx9VfAbGjxAgEgLxY2fV3Afg5yhKXJ8Xfwfc4T7fLIrMpzIRtAU2WtB3cLcl
kdoDp2Od2iZOI1FfpRGGjhz4Ymoi8hX+TnhLDMcLStjx8B2kvwy4WXBWxl/YixDaFPVTt6vDg9ls
Afz9n/GUMa6/xLMTeGC6mE75Yea0n6UIuuWqMujoyafSrisIm32/EPVPmjqewGuCD6NWFdNofh6D
N2C0aiOUApgsLZSGgEKHX2z1uFgEh7hip2pRoRuIURl3tTA91VOxix6TFEMBWPl0OPal92J17K1c
4cU6O7nKPLNb7ItR7qJiPrzfcdFSrTNbLWdCx2wYFrx+YO1OxjhqXG25qZamx8AWTcrujfKnsGu0
5kaGrrNeB39PqzsUQBSkpypDNatA2x3hbB7KhW34H39GvB7jJg6wwpDe//I1Gfwtsi7CkqQVmTif
uODvqgvJ1MD1gOJg0jT3eI+rwEhXNGaNCGOTeyLSiFLrMfUAbMuxoD5GAWOcBA3xMaV1v65x0UWC
b0ydab1OdDyvbEy7GW06zqscOPhxIDmjxZzKVcu77cV4NoHtQdXG5Mw+yULLoGsA5F6q8OSe/Kl1
p0V6CwB5oQ0MXb275bVUilvTWEENctJ1pUgSVZ5c3ziCfaeGhBfogxUYtTvYIjcgHAUTjzx5OBzJ
ECQAtmfpVjsVZl1jedNF0SD20bSOgTuBMXE2jNUOYUxJOiVGqWrnv/KrrNzBsM3uCpCcffqtkzc1
Ei7hJv1Q6zfAhNHkZXeMjzceHZWL6kR7gH2iwjWCnHqyVu9qXQhdgXzAFhMQ0rCg1+k0TmP3yFYE
kRgHnyTW5WI61RI8I7x+UHXQGsuQRXNa8k1wpt0eBxkKGiumenkbb9epbHhPqQnnAX9R7abyd9SR
bbnjR9p/oc66Z6edxKJKoDqLusPNttYTFNo8FsNZ5f56md7+Twbysh0B0XhJS4VLUYfmKuZq+WB/
7rGrrUAGzNnHYz3Dl5otRedWABl00M0q6e9l3hX0CBR9xTin1DxFPYC97hSaYj0fOPFRkcskgNBV
Li7igqgeUxc9tJPPi/pF+YMhiVUtWIlrV26vXmOLvs429KGEgQnks1m3ySbIyXHMJLq0MPw4hSaD
4Vy3QJJpbK6k1lEEUKoGn/jMN4z2mingXQB12rmWNjAkrRpaX9j3cObFG6cPbYp4WrLcqhUy5bj0
GSQtGaVrZZoQet8trRrJ20RRITVK7rkR5W886pqsFmIRdm/PJi2mDsgjQgoOb+Fxn9kqZXXANsZe
ecIDAQyZGnYdzu06pzfEdanx2leCXveOb1xOfaHF3Pw5tfhl0udfUzsmEn+tVbMYNJapokqYK+cF
EMLsd2iEKm4JXatKIPCFaMJWLmKTII2VSZYZBkHyD/VuW0RO9R8yR1OirpNrmGRrM0lGp7b0Ze9J
biFW6GMwI6RM+4Lp8nzGXC/nm6Azq7YxdwCzv2HWiap7vPJirBCZPw/36qe7Bx8fFviLAl5vhpwR
kwzntGWRxmXgK7Xav0NZL9SzqOINQEb0Eodv9WOQGNdI1LEJQLxRIBAsu1HAIUlhPqyHdiCQ91hD
pIfY4iH8yVv/ET7Q1kZGThDBy6UzGbLyu+r0nAQpyzTJSb6hLAbTwFUKwdc5f63gd09xGhHqBtlq
JbYZ6EwyyNacGWRkARocGcoB1HfOsaW0IFixtjw2tYHG3JX8tdrRm+zW8bEXbrMGxuPSjp2Oh1tP
6rNyX7OJRlDP8ZxPSHlHxUo+PQHNnPbDHLPpfTQiU2jeX5Vk414HKxS12LyBDQvD2HmooG0s3ZKI
KclOtQdglZ6goTTAoR5vyvFyz81BsHx9ZItUNs64+2dcryXbSrqbiWe1klupZvA8tEYBDGsdscHJ
RPDrYqe2vq+bCe+h1xJIo5pr4xPcmZAas4Bd6g9CkGSwfJYDa+j/wGGUglmxoIVxnlPiANQpdxaz
He+TdfioNS4sKoBCMnqcAL9tKsa2gitUytXgrTAdOqD7SB16eM8UpY83fBunjm4XToIM/Sk7GpAe
vYvnQfb0S3o4mOc1MdAjQ8QK2wVQoe2LaJl1yk32CFj/eouQz9TzQZcPO8yLK7jro5tpZsLzGlaF
Muu5nVAo0lVnLgOKfLx+4oXKFm67z2YOtLfCIwCAaZWLhMiCsOB/gW2p9k/BiznXT+8O/dWHnRUn
QauZdIregXv9Bf3n3hMQIT3wrBEdyBGYP80NQENCxTyiRpbTUPMkpICJqxYjKX36iEWGVeMcRuHP
iM2I3aiVTLsfPDoOIZBUd1cyXfs57n+z8Vp9AAqsgBl+JS7XZPrCzBmcsUAKM+Z/32b+Kjl3F/QT
ipfZ3dBlr6wF9bxsdJeIQZUTwnadjzlMl2VaINAdF7yVSZRxys64w6Wfr6FDJJhZoX263TdJPtcl
VDTpH1BNQQ4YGlWynPJgtLzIyXXJEYeLODVoEOSfinMTWdht0h//44qQCy6gV6NRSQengehIwuPt
9Xp3IECvEZ1jZYRTnxZ/stQckqQFnsZYp7tteFGJdsJ8YuhFFw8VFeX4iKrDqIKRfFjn2SC8jBIX
7VUJpUS/7zJD5uC1EIXEn71WJU4u/LncvXz+KsqP6ROJLdq6P8kDvtDMJWKXn15774w360/fRsgD
EIyQ5SfrL1XF/VTdFPd32IYNzSMCYnfYyuFPmG+udKGc49s67EGJELW5FKdLxnMpSKHh7d0SeCmG
iPBDz91iuzWWFzMh0YQQSqfkLrJdF5JK27vubEtPBAeEF06IhGC3jj/DIIPuslLORUSj8yu19Bbb
3Npbf95gVVns4m+eWvuSCRJ/6gtv76thPQkm1MHiRU+cIFKO459MpeVqH68fyN2TnoD8B31ahThk
s8Ijc+A3ugnr8V/LMbb9sqRqzkIX70g3jQBwvLeQisR/CV4YngXWwwjcZEjfzi3Y9iDNg0NXwJDQ
US8/J2W1TjD9GG2iEOrX5iskSfM2pMoYZz45Oe1NmoyLWY7XhU8VvTtbfO7hDi2NYEtvXVGT+w+p
eZbuWULNMwUfLesamrCSGXQHT7pYMfbijlPsusX8saSItOTIFgCaggEqoBXRkbG/eBqU5RTFdW/o
dVFokMOCwklkYSp47a9ND+vge+8lidLWIygj/TpdTjaYekZcVsV6WJ3GOmwjvia5KIOnN/3QSMIF
tvg89ljLoplA0dJnGrP8HyW53zhl3rz2+5aOgPv5KTU5NQoKvX7/2vkoEhhIBcJMS8JX7gyHcZSw
FXlmLYPe9wgh8iz7IMdElzm4cgh+/GMbJXbhkyPu3psCKOce7o3w1lbL9ndZctwKDdCqwqmuKqMf
jpnlp0SR1YySCZew7gJJMIghRvzQRff7o5z7cyEpQrjC2r0Cxahd0u+PwVl4sLNUeP2QiIZn29bE
iCpxwBz2R6/OhD0WyX58l7CEtpZgrjh9XhrgHC8Ojo7FaYnwlvktpjA3zhb3UlbJzRSEhxvOmM2M
jHjpVZT1vm2SggkqtG7TG29PDTzHphKsz5hwWp9c4DrhY+FCg5RcASdNesXoFN2LeDpEFArAa6ls
cwRH/8bGKJiC5MB0QnvJvF+CCfMvc4DcmEXb71P93L+jPXHwBZh94biTMs+97wNio3+oTfnEw2LZ
3xogYSb+Xywj6jaaIQkHPrdEMXChlYXuOiE07tQBH5YLq/XeXDhe39DdYwRVfQRO63FqsuoNQ55U
4XwAhdakVylxg5BuE9QUopwj7LeJGRnovFOisT3nGU8AAKPWArRe6sHL5yaHBoLIxF0MJlo8OgPZ
cogBhRWCXF8W1k6wgvplHurd2qGQhlSGHkViYUVICFximoTGwd6qe5Xh9/1CIsFtv4/p4vQ7tAgN
7GAdhyzTTJQBLypEO6OoDg90M1v+CLUH29OGuZ8Op7+BCM3msMOUHrceQWCZvNSlabJe3ggP7BvR
2KAmvHl7RQr41Gh0nWomfOq0uFnYMYsCDdym1KzhRINUSSjBNOIqBSzkGJ+enItWA3ByaORAcRYG
ecmej0uYAdHYQpgpqcKvplSaBe872eaiz5HgtEi73rUzey690VIU5+p/RXZk04gnTvvBDkHCWMm0
xaYwBLh1EtDUih0BA9V4Iwr7fEW4kUSD4vapGUSloQONsWvzFyAhjYKbmS7TaQW6eyUNby7gfIpv
G1jkbenj71EYoqaGc8SOXIDoM3pdszpwH5XEEupMpDxmr1FecjQTdQ2dJJoHn7xqVtACO5ELClpu
8ye3/6ZTKpKFxtfJbc6yrlvWoGvljMjj8yJ6TU5vehB+cHSEsCnEHOYnKYmyB+AKldkOIc2kd4Ig
9lUFfBo0a+VUUVceBlJ5SUwiJw1k3rRJKVsVQLro/Ci3yVFDFyV3dQh1LZgV9kEYTurE+iv7E+gw
rMPXb9nvWYJS9TV0JHItE0JFnQIQHdl3uYiiO5B8OccYb8+bxySkp9VddgLvR0ztc8kqxoVGXZ9A
a7Fm2FSTEeJcmiIYMeFbrebyeY53njZR/VKyFkk3RVEqjC9bfcyU5SAiR36ksKT7m6OxX/WIfT4p
vmF5ChIfiKIeOj8k9KMjgxbY9UR8vN3J3MswhGbtuZKuWliJv0fEoM6j8ARcIp+NtUJWEYRNVq6U
q8hLe9BIn9eMhky1RqeVdocyOguiy7Q9n8HKgbbS3CW8GKrVowQ5HDdTuRmEkLIpAtbz5bdlFVYH
IQi//WEAdo38p5d2sdZBbeHwt2vDfXYas6eu1mt/GlKVJn48PPP2YN8OAgTjKDp/GPUj5eDPn/m6
5pJlTD1EMo2bKQ+xVIrnDEYKaNDVAzpwCNoBeYtwkB1QlHq8amSTroUk6QWFfItN7WCj/l8vy3H2
z8WAQsIuoJCW/tt+TCcYGYEXuuYAXkoGxQ6F6tUrgDFtyDbMNze3X5ZMpAPReOHLRURbMn3eizHZ
prM+/up+CgJzf+9oTW+R0dUiKoh4GFOjWCT4AfEYVstl1zWfilUSsNIaCkQes/JW5OMvBOu8Jsdk
I5Ao9bbpljOhODNDztZIY0xO8BDcpnoTqGQqhE7G3Ev5qW63Pb6X5kYEEbHi+tghwsYYz2u02Yc+
ziPBeVfV7ZbVBL1HdUynR9hxs5ErcShM+rQrIv77TELW2n8dgbGIS7DN/MkNZrE/Pa8EVeIbvmbK
EK8T374jMRLROYzd9LcqcUvTKhi5oO/lyhxrUU1rEcB7lmCKSXR6Mem049wsvyFvuuUULKu4szEk
46a1BZXHtx/reanH5b6dMQV8lopHdhkTOsL7ntFhkdCqCIjfnV1b3j3hNLoBXiopmof7+ch0zrCi
2MajY9aypPDWYnTOfQTImpKy2W8NnbONNze5CCps/mSvyGd7eji99CFaSjsj41Xl6MaDDLbsSQUJ
3NdX1auP8WTAPU3lhDOaVTc5hXKflnz8WUTEXM95Hw9pwwwNiqi+FB5sYTA3fTSQ5qHjKQKswRIz
rIxtAp7gsfCjqL+UqLJ4L+qeWUnXt4zSPLJqc9xOjtstXlJmLUzXjuLFdgDmKRTDZCjI7bRUGlUc
K0DNxT6bXGeXUn6+W7Ni7H6K/7kb3K2h3kICtDGmFyVpMu2JDAt8OYV6uXTxvVBDRmYhf6F1lNg9
DRNuB2+jfYuBHrEr2UE4rPLflfrE2xPkDvPeJVYXoR0iekf0AYk2wLUdwDa9tT66wgf13r4n4EKd
MAx0JeCcLX1oLuZGg6uJwmDXym5MWVk9+zIP2lRQT5QU3lnJCY+95Brsa6ih3K7Qvuuju58hll+W
pzwknYjOvdhlzYX3Rn2WCtJbWqVFK9iYtmlut3E6LZxbjAuQSkV8g1kCPN4SYQVK7wjbJT5A7Ban
pPITlwqMVt/gQi8I20G/cPyDIFSUqQUA2QsKnLiK8+ycfE0QPT5kx7NWNSqvtAo2NiyvBUDCVPny
XUEz8oL6umzldXe30bsTjMURsE59416ax6O40RbhA58R9fXwH66mRVL7U2D8Lm0p0FiNlkoHL+S2
7/+yZfoRWjkN9oPb7k2ePYsC8cdoTykfiODcQojzk8zgXwKUY1lyNS5tlCizWK+lzSzJayKaQ3Co
95qlA4FouoLApynLDYPopqIepshL6ydnoXR/IGaMD/1k0feBRaJJ4Oy33awenEPRxs1ZaYksVGza
GcenpAARvtsLyXuv5SJ341JNewQhuuiTA66XHE62Y10z9DXktBdKAjt0Zk3f56T2ovvdvXELJCXc
Swhwr0baoMVbIaax1WUoShFuAZ9HQwkqjKbh4Pqo4wvsijT/z/mpDGvADFo37NbFfM4k1pHN11Lj
IytawWWhX/sgaaHsgsXv9Xrq00RAoa0qjeXLXZV9MLYJlmFQMho3GMzCuMuoSGyK2NiTPsP75ziU
BwJIRTpAhi0GLrxlzvrEOXGDVdrmjqDhW37XRK3tLaXtxqPPNcUggFaplCAnjAKfihlRuD8GSNNu
44gIv0Ic3hMJte3ae41zJ8UQgIUYwrTMeTwfayfuYcHPtJV/MBklCqhB+zfOc96U8K8jc5FhqgMR
f2K4T/o8IN1RNPhV7K5u4W08OAnQdyoUks4YfRBRq9ClAgt+HcuZbD5JSNJQnGzl7lW5b4YBgKnF
19vP5JjgygIFDZ2B1+fM0QRwum7sp+TN+aK3/l2dyRGyYQ/8RsaNqzofSQP8TcU6D8WgncGv11PO
MPn2+1Wp5D6aK+qbxhGIfBey+jmiGAi45T323U1xtfGlQaZLbv6J3RQU206+bYgsxiC6vVLBqI6S
SXjtHUIltimp5wBBdtrIniwRfzEtX/V9tOns79Tw4kg5/B26OYjSbY/UToqud5wiN+qbUfz4xCPs
RPZv5OMC5S8zgQ0MdiRxiF0vpQ1Z6YdtIDs947C2OpsWeMEMoI3BP3AtUiRdEpUGtnZIVOR8Y63M
RH5t3f8Rr4qQimYMfxFlIoeS2gquIMc9uk1ivzrBh2MAWaXPGBTdWqMoXrX2iWjCuENj2GmSh3BM
nUwqWFeRvaP7oXwKGgFdNNm8kGp6bBp8GqRI8AG+JEtaDjn7zEW/hHguC8h0tBwX5pjhNTd/8KRI
odu4ctFDYT6lD4rmLBeYax2qL2BrSDydbDAAou3A54rtBtI0l5qz9ANHBrnDB5hv7zocDhXb1x9v
sSECuSP/lYRbGKb9C9HqHobpq/F0Gwjk42Il550rwbsTax7iR/MXgmlB8gm3Tos9ydsLgp3rpj2K
ym7gaSC//gT35hZ9ESIbRLPZlHr6mApypC9I2Us4Ln3vyyptqsM91ie8gFjdHq4axqOSQH3OxHWA
SWF39OopkUMPxJGTdpqScNClHfbAbgkX90r3lt+lpJjlPFo+FMzCgVvzzyS0LgsA/RtUAM8z0KZz
IjX54sNoPLcRpHnewmu3DQW2RWEHNhVUL+61gIaeU1Of1zCOF2v7qc7drQPrC0bhqhuD1DE0tZgF
o6IEoLNRv/Lm7m5xxAPvLfaw0M0VWdaVdqq8Kna5+s32Q8ZYAppHg/UTTKpY7jTeBllZvZ7nZkoq
6nrLzLQIjRwRmbZmwNaXlDktYE/bznyqKxF/xaWCf7LJ3IUQLIhddkQGWLsQeIaABuwkZjhLP4Gw
SigNSdl1QlcFDyFfO4Qpw4TKf+WD/mU2T/hXyyIXLZ07W1mxisikd6GwAKpmSWYQfCP0SI2cN9OE
tdJ7LEVpYfTmHJxEPHmuL8V6gDdCJCWECE7u5L/CPIDXWkXLF4g6fKrurPmoaH8WxRmzz8OX2uIT
VebWRy5BTOkY5G0KT4KMR64aV5KTl0CODkuiQwhSiDaMe3FnwLgH3Ox78FNGR7JrDcYvCw1x9/mz
LkUX4rnzA70za5S6RpfaIl01nKHR6Ck7G/llT6Jp5wq7ikyOVrmKkLM1kclKRL0Y3hKP6/V7Qi2m
VXOiQsJdoFHwf2chObUJsmoYBcasLtDT+Ukowi71bd00tZz+l9RY+q2TdUpMUsqDd3ohVUtKoDng
Act4az0aIOM6ltqkj/vowEetjFco5sbRGNsbbiFvrwFqj6M6FYnrKSlHUp/P8YFBcFJmvXcUFq4D
hB4NUv+PVwvIwnYQkg7LKwgc23SUN+43z2JtwmeFx9PegZPScW6vbjwLVILxu24w3rGciGcuh93t
3yvHnnmxMqAi85VAe4prbVl6uoH3TFZiGdBthiIDOkSlqxGbFSU9KwLiHWid//4h0ryBHEDsDblQ
P3yFbfm7DAaYQlL91KVfjF9ocACR32J1PrOxa7Vxcd2fd1FI1x7DDRtsD607XkXi048Ln08SFWor
kpmovg+PHZ8elhOlvQqPdd42+Wn6Y7PmMaIVXL1IcBsBMi7yeUSbVOKMcP5jovWp/w8MYHTmKVdR
wwcrjo2U389qEArKVxTtJAnZn+6orbs3nBpaXzfDB9ISKFG6eYTJS4vHc5GJD5RdU3YBWsVX1pWJ
lnPlMn2fIFJCk0e1Fhy5Rna3vhUxENduk/ZmcXUeaqcv4uwp4amw6jnzHEMABN9/jXV9z5Q5Yv44
BaAHhWndaT8KPrJssxjXkKxHe08iZjEhdJlvBFvAuVEw+Ldkjk30uyn5V5pw7XXSxb/KNoku+2Bs
levdbOZGIplv77zGDacxZGhCjWKbzj+51TSdT6cn/ZjHzfSOWpu33+rqLRu8pT2Y+lQcOYisgo2H
jRFYRzgESF2hA5dA0D1Wejl/kovindDkfX4t00cq65ffbcnUBHW87wyFGY8WK561RsFnHSSTESv1
viTgGiTMbpJJE9ZEIjhSFyLl87cUE0WuAnsfOxgaYaNuGjhuePhmDpp7uDr+BlxWq5zLKbZQev6I
SoWNmiPsbDLzkAg3le6VCR2UcbVgBz1kJ/4THmMrbjvVV65AAc3fzLe3pRSzcKbSWaZQDRRczpng
Bzc+hluDWm+Ez1tRdpewGkQTkCFSNH4rJ9Lc0PUUhh+04JSksOj70B5PXMH8u74UaqRuZXoG17yf
0db77Ndi/wW7FSnl6FO9zvsBTufb/0mIMPk+yB1XGWXSsn44YFcvMJ0u/zKlKuozxzDkAvptZBVh
rLtfCoMGV/Wj2mLP0J3Eezca+8hhDMudvmHH8nRHhUUhztSHgKRB0ezvCNbLE/PUOPPnrRqvBPFr
0l1Q3WuZa2eraOgYvae1pt4uc+0BbYcw/BqISbRbskmLqXXsUXh7dgmNUGLnMpY1IYXAI7uw9oic
TJF4PCmspHtgNw2QN+pdN7fVlI71rT2ugS3kJbPttloD2F1gQxgWy7qw/cmXSjXHyHiQ8KST7vig
0grRahCIvzZ60IvphOe4TVMtNzTOFRjypsIR33ySAFihwwEhIM2DQpfVJ+kZM1ncPsBedBAjPlFe
jfXXsDCAbqhwcGSbW/lvj+R+lASXuQYZgCWjLJncnvnfqy85H9I/2NOQ4pRBrj6KjfmgwEKJ3N/9
RKo4R3qdqUWaY/JCUS5wMkB1VJNgCeCpwd0TUoJRp0rPwvpCp+PIs9YQnxyZXYM3I39WP4S84jTw
ke/SMvq2JSyfUoOH56fHzdP2dZAjD4Ijmwpaas02C1THzXIzrxZPtoy3ryX4m2xSjDbXOqry3m99
Ltg4YKTMExuKAsKN4G/UsarWtEuSbYlevRnLQszqJ3pp9G96xR8WyoWYuhFLg/A0zh8kcujh8/QM
m4VirkJfIJMkOVWhl7ugcWJJu2A/g7EOgEZqQd1txeHGW6FnjlWAvwW997WtGsU/xJpw3HbxPUHW
5Wc335UQE22YRpCy3e4jLSgpPX93wo3Mdx4LH6ftdjlmXUat2dAC9FSUx6n6Vhy5qWw7YmTyu2ER
cidpVRLVXI80XHGjT2FQVMqFZTjS44HA1ci1nG/dOcIx2poVNOvarWv8mNE7Y9eo3vgiu1MNS15J
zE9XBE3FNKQMkLRFkNckrgdTUDGt0xScydHID+zBTf6lbhR6+TSvWo5Dor5YJwTYM89ymTxTz/cz
VMH5FeyJDSF0ZJ8s4nltHEHKMqoPnuNdfGfnDsuf4fvV4+EfHMxtVMBVHpFyk6LTzXezrrlLUX4m
chFy8BtNAaHer+ZaX1ue6mTpUyal1kjtIjhs1SBVccRIJ/Ur7oSd7tYLAI4JpOcN/hIbeZXyAXQt
j8l3+UifUfgnCo/qTPB3U/IU4L+rWRBT1W6PSpZZyC5kL8hsCGoV8s+bMMO9XtsbsLP6d5fKaGAr
t6eIvJvznmoWM3inB9/qcUqMPkm4vJIzBzvvQ/TO9dQ0pMvmTWnKQYhYOWRCiLvYoPgKpWVYwKdo
ZJF0k+k0lXUwtJuI49JWi8M6haYSPl8yuyE8R2f2dKb0gdbd1dJ9OEnL7qICY4Te/Wo0jdCnVdof
6/NqM57yBGDvdi5YQxcedqUCknjlB1b2EIcBG5W/R/gOx4YpVZmRguywvtjRHtJMSoc2h+yj9+2U
cMhJmMwqZ0CqgKKIR3abdVC8V4Un/V+jZBr2YgWvwYFVnUDfviaF1yNXIqXrdEBQhFsBjalCDLIi
riUi8OUqpPy7Cp29UU59NAJBhAQM31sZ1Lu3Sf8OX+RLwneiO/weB4NHjkfafuyD2rEfT1fl6TcT
H2q4v32biprwKCvY+KU1Tej8GKbTimZXqkSacyFRUkwQhS27/iF22g9JT0KNbdf6JfU83G2DlWMp
5Xlx46R4+7XOUC6MqYlHhHhNSc/DmD/FWRLrq2f/nFbFbWAMJBd3iHYU21ax6oTFj2Zr34L4aXuT
4eRYTDvobuQhOPJUNjbcdAY8bU2IVCjEgsnZlHwLkwVTGHm67jsMMHmmeCm6taAokBaGEOlUIdAf
xsbwZU/J3jQ/4N2l1k/MQdfj+WNlhaXV21SEPDfTN5YlG+JYPZ2d0ukHkZTC//bi8cl3BOzAGjCC
wAH0LhCMmgk+Iuh1DbRjiDgOxu0ukjUXglNvZpoBTTZahdboUF/53VAmFrEeI7uyN3SZIk4EDWon
a4KtugbEMDXDKaz+4i6acs7VxOmiyfa/cbD1MS3wNNo6rK8QKQM7drncDVy2chxTGDcSuAgjwJua
uL6rlPXhme8bOCNaJ5k8727PjikYKfbwq7BxiCsWrgmZLPpnW2ksPCJSCtoT0wKE9tQY/onAH/zx
lvifFLEonUhFqxD7Yh/XAcuSdnSPnm1GtB5cgxpHXyUNEb3ws+8OSmEWY6+oOsQcZtMOPxQWuLoH
lOwTy66GeC5npJuMRN7dWfgT3/G4QdIW+/YUR8SV4yw0zV6r6T46T9TWBFqLRrh+I+ADPDRclERK
GAb6pxd2tDZfvY89TBS8vAvxFl8GesbBicBnODU8BkoneNPmv7IO23ickisUbQrlpoc1DYdD0gz5
mlKmc0DxFgXW3LkLWMMHy5OLK8vsAt6I0QCaEUSDT03EjxHkVvOYPX7EsBivWsJj5JS9t/vWzkvX
74s8w3FPLscUuTlsMmUxQJ55wM2OIOtNpyxHH3HJSHxF4Lx1YnnCA6gelfPsMm7lOPj6lHNOYXIl
QEY1050bV4SdWyMvxT8HhuyG3z23MmKWV6UvVyGaSCVmkBMa3r3RSdnrlmh6Li3N/vLlppWb7ZEu
cbZOcSiVe3HvzNLFeSpinzZnaZBjGqQOeIxYwl+Sr8YKGYw7Tm0REgaIbJ+SZmdBArG8YpygtX7v
FpZ28muizZ3beeTM+c9QN/QF4/rWRaDrVuFLzieb6m4rUVwWcMJSE84V+MLxsMDkVKIDPoy24CwZ
0ruGCovEs4mtjjQuPOWxQtUucow6yyoDpMZ+L19DHBIan4bVnaOVwYdh2sz+WA0nA5uMReN+PKIk
cT9SUayds7wLwoRJmCtS5iIvcDYJpG63+kfOVG9OE0khvac8kHw8bMLRVjHNbQ00HSgGTBjTYltM
eBeOiTNwa4GKsKF+7TCHRh+u9ICBnNKB92ZsgppYl53lR2L/Gpv9cjKn9sClA2iPlhYPponZkaTu
EG7DFy9tAvNFw6kwS4W0LWSjcMxHThlFY74tifk2N92vAAIJ2wL1LekQc/8J8PVIE1s4WMCsEkFR
/d8tWiX1b5856LJ8b6dKOnI9Hni9wLHqXgFnqikEfhqImDJrXowGiUpExcAQUFUxhSAP9PygNGk5
fGsTqT4vmpa0YbbNVV0SUmA90yuPakDUKmN3fr6/JLxx9SAUuxQSXk03wd0LF8wJHQDgPxYuNUJw
SbyObn3gXzFEuG9UwxD6Qo0AHZr1nO/C2DhEV0VYMlcPro9n2GRV1q8VvXjORQ8MidkFd5WWxcvY
T+C2rmeuPkxBlYkLgZgA/pv/oCsd6pc7z47CLNXnXpCo7voprQRPCbM+xu54FgxV205HOOzOBMeb
NMocE+LazyHfTrGUs+Sj5RIMqTPoEORAOSW/nKko1RxSgNxYWfAOhfoTgOIwCId3jm/LpZ1T9lxl
cnuBXsssDx6Qc3X9NlQ804YQbqLtHFOd3Z9z1kds7iy7uzD4rNpRNRoUnG8oxUqZxGK7rj22kT6e
8CUAJeqHF43rFAB6L31ALEcTQJT/wbXlV5vXouAypzyYuJoz+N+a8dOCrQakNKSNLtf+XAHxwLSz
KpVhLXt5Hkbaxqjbi3zG89dSMQTc0R4uSJ2bXPv/R0216M2OO/uEvoIsIqoMl1SEQ1QFwbWp6D1y
Ashb7fWBs3CeVRIKOZod3oyteml7fQbwwh9Bp0HzgCR65IMY4p+xuKmVTaOszMBuypw8PeMbRcdd
pY1wCDQvmyj14Hqas0xoDl3ONyPBAk9yIcQ4PmZOWcphalJ4zYr5hg2VlRwxcJtI9/V1vtbPuAXb
SWybMCh/vWrqqUgVBPHoFbipbSf/l/yEuBnfdlaOTKge5v8jz2JO5IIcJEitiTGcL+UjljZfulWg
Vu+mQysdI8fNIvxwdbu9F4fmBrw1H99UEtoPd3BJzNVdFMYiH+U9DkVQnw4LA36E4cDDH/tcMM7g
30NrNXJHOihOzcEqmK4J7OVLZh+Bf6vwWzKEwDUcfrt668tFvPdrYyovCa3DgTSqNsE3elrGicj0
BRygCrpFDW6noEstCpYmuIyYUgaIH00uYaRf5SYM37JfmrDaZdZmK+BC2kWQ7aSOw1W2Q4ifQkBD
Hdx1vvNzAXfFQ9h0RNykio+AGNvRnWXZCVWee4mdCMfJW4QX66lsti6Y7H/Ittsaf30w5JaF7V29
fe6OIwD/qDv2K3P1owx6h2sXr5Dz0q5MxECjA4bW4dIJsTqlZaj2UOGg3tvpGIv3Xyh0xNncBTpO
LZ08LGSBxnG6wXXSmUOrwKJOU/4CLMc8O5NLQcuXCf1+TT34L+kZy242XJ8hUrG/Ew4XqEcx2ffY
Z2Pir+7JNXKHOj7q/ofBPN0pQZUEeGg8FBU29Ejmmj4YjqlXPCNDrbIh37/F7PN6EIxS98NWxw8Y
3Y1X5lD7HO95Z5I/czqldy4aY93My/rdiCSmN0bLF+MaNIGh4E7b2N3vVc7EPZA4iiUel6tfg8QV
ihdAabdV+Dd4nLdy6RquwMwcrgGl607gTDcp6/tyM0cB2YdjTtXBjSWI72EedGzmCFzSO+DRR+es
ZEAUPym6yJ2lBH0a8INMURVKu8jM8agps3F/u4FNJ/M56TuIOWZikeFvIBsCe/G8APr/hOM1S9C6
RPW/+TwACcX3a7/BVzG/61yJAqXyLCXGkir+HDuTXOJSqIcJ7alG0zYiLYWN1FlU6g1EC6d1JXrh
ArkohroqOfVim/jUXVyfwEriIVdm3YA56YWpg9mRtBPX98HypAOgXaZBmOf91w7lBTQF6/JBrfdF
EnX9hlUWdRBeApvTY1qKlR8RTk922M2JGHdn0vLCxlRWhaJP5uPBES9kpBB/8YmQrV6Axq0ltrkr
e9a4bqrxQv6+gmApFL5CFpl39z8vX1Zh0FS1LiGGZ5MBqNq/lyXpHn8eQQOx14UYeqnQLXy2MQYf
yZQmgqlBWTPIqg+p83fTb/AESDLzJCEhBBeqzgJKXZD5xzuhYk5aMgU6qaTgBnuDgCuJh0v0HMn4
fSw0SKD4LrZfFucHlpBWWo/RsnoGBWEBVq5gMr6QU3mFEcn6cgpR2GarGPJZMCtqoUqrMcrnlF6T
DQG+LrsdCcCVTMp4cw83QnEzWeG7AZ/FXFTO0sptlKuJTRsPUZM5aIWhCxfH37b/exVcpd7fC+xh
+jnhnXlz5D4xgPSGcP4n66owJ6J5eJc01Vdn/BwvOXpDjCh3+qz+veWJCaa3HrYoVpWxRLKdveUh
/L8fm9YRdSYhq0IQgbeOZYS49cvYsMURAa0uHIaYsF9tOMq9Bw5ZGqyhGpaiDYitrjJpQapLrhIu
+2pqI/oJXnqJUDz+F7ygEhe76qlLVkQbYYYJe9w+tJKJOEt1l2KSllQY/wMZ3e7uWrUr7nQRXJ52
JVT7aBCpaRXJpyPM7atKxBdtou7jyE3or9cpRmS1Sn5awIyUO6bFgAw6XIfFTiBv3E/3rB5RDC3F
V7IleoV1ryR2NoOdklnpHu42JhpeRKrvYoIu1H7wm+1U3AOMaiPOlgKA/62qHImXvNEkx3vv94AK
0X03GeyBj8+15RwhMjRK5/vLTaBSq/VjYXpUnBsfntijcf4iEGkQXpqPlmGi0CKPTy3HKr06I19O
nRXVVtOAeKCznZSA9/EHVAqvV6zyWAlnUX+kYT4E5l7OaCdWzvYAmJKEBte+bnXK7EBOXDTRrdH9
C4E4T3l6/HXoLFb0x1Izn2pSA67T0J06kjO5KbiN8XS6CPBqoUJqXY5sFIJ8Uc58Xncv7PopQZb4
DrxOVKGWH219dg4lpeX8rv16wLNtcyAvG5rfuVo9QWKw1GWSSdMG0lPsRR+LNRl0/QnTL9bN1Gyb
9XvLnhgDu9y8aCeZMwpDcoM9M8D6Fthjc6cRk0lZiZGzMNGVb9WbHNhHUcN0wsLUtpo5woVJ4wE0
zzOlGZslcyP8oY2OOl+wBD/GCZGCxEEHOlxUQlWCm6hUajVKrNPgt+fnuKZ/VIFRaJkvLOw0osHT
8lI7Nmg91ujoREt/uGGFwL26v50fxg9bW/cFZWs5TCYIagLqbK2WCpB6AEvTtpTcWAauabxxp281
itJvItO2kziZJiQf4a7w9E2trosen/q1RvL904HsMy/pliMBoljWrLh+1EFnHzxehMShy52D0pNQ
OthC5jqQmEg3wIJgl8Y4EqRE3DIMg4SHDunPNAKfxUj9h3xaP4ykZVWtN5vKzi3LDJ7EXhwHje3/
Cbozqc6pcL/+l7Xu4v7KDj6BeyKHpWiXNF/dCt+Q58mgEsHbs+UeKG0EHAFHOLxH9IZq8sUanxWv
NsB744Ed9FujbbtqnF+t9sHMsFYbG1ffUizWsf9ztrWNQdPbJn9Yh4oKlkMj7ZzeLFI+M2w9WYRc
PRlI9CYvG8mw9l/+PKDISdmVkRv8Gv/zvZZJd9vQM03z5q+f5YTPaj15jtFuIxdl5MYyuKGoNkxA
mssJLe7jIuWdYiXuT8FlG0Du91bH6qriojjwWOlOIxyHq1WvxqzmuHLIP8kYTHfZk9hT7xglhjey
F5hZ+QgCxy99yimAuxh/VPqE6hcyKvxjoQ8cTr8k36/I7uFuAZetGKValQReKcCA8dYb43Nw+uHo
puKDKwRurK+LFsU/1yRcbiu4opdV6fs8EU0N/OiZsrv1Pk+NTJDs1IhtWWHebcyjSMGIDjw1NnuN
hXDz47rDXYEm+3cQjOD2OFLlW+h53oUAsbIWEW11r/tFgxah0iJhljcXqiKnniRHDcBgduYiT7Eb
TGCFFVkYpXtokU2vMnTwEDFA7L49M6se/p71jW8YBSlBeojU8C/Gf5XSA2MHAf5P9jGH1PmBm8mi
sbpSqEk0Iv45alE6Et7Xw1r2H29mtK0iweEqD6aGG9hGHyW7WBHIUqhJ/pYOKA3lVbbS8W8ubnZ5
I08ucfSJo9vM5gXCnNVtsESBCGVhmA7sY078Xa6X4Di957lWfZpOaA2L6ETbvx0xojyxqy7pf+Zr
BgyId1Mmvb73/jqjqWAQEH9H3vigOMHUaGP06kh9hDmMIIHe26mISi1aDGx2TEf31OfgksCRHHG4
Djo9rigYwk92qiRV1nIbdEm1+BS8curUz+alG+9ySsLi90NYFYSVjADDUzaxCGMRGzJ/MtL8+xp7
pIkt1MuyK9uiyf8aTn7di/ottNyAiPFEvFPqa1EwvATxm/B6huZrF1A9LhAE2bPuea3yOW1DkTgF
Bu8mApQHg4UV2+WxDxKZTJa8nfs05BmsqtBMSKTCx/W2wsN7gYtEX9hp2hNAgFw0EeUhz9TBCPLY
sKxh2VKot/vesZUAXqbfOL7L+c9N1MVNwzjwLTNLawojnolsMYc2M8tyMpJQr2PgV+J5hzzhFTD3
cDkG/Se+bnOrFxda7lIE9eitBlZ6Y+HCT0ooXKmbh4oMmzlbdqmikhQepbc9u39LqRK2PdniZEqk
fypjWrH0icGme8wZdjfYxOsc5lxXzHgFoROrkZ5+21dmC/GqTPNqbN7fqfvVpWejUPcnhrYpyBwL
/E5DkuriCCFyiv9O1LvYtlZJ+Fm8TPTLjbLHi4BdI/3FDVXeREBbnmEu9OtJgpKXzbyUMZrcBf89
ASA11tYlfPjaKQtCABD2j1v7kbTDCOvXPXhqy1Ji8k/FXw2aC3hmUbtC9Epe9dL9tab3e+QAUbYE
lek1szJXzXyTbEOmR19JI0oWYgFO/EVhJjclFuh16Q30JVmDpzYMDv7ZWRr+hEXSl6t5pVCmlvb9
ZMn6fUH3f1z5C5YyJ+P1TBWD3U1k5cunbg32+pwFknIaDMOQuCtr7SfSlzP2z+vYa0Hj4VGaHqXn
PxhGdaTnqufMmVVPxSZTX9wtVHjMufpdrkLuhEs8amP9d6A0Zf+Jr7hBVY7A/r2nL8uS8mMhfEq3
CKpM/cD5/1zQk6znY2Ysn+Radd/AGQe4/5nbB2wzk6hxdgIiRZWMr3+A2OZEySLIgkBmZLTI/Whc
8D7fitB227grBuXEXKxdw9b09dICyHrL3YcD0xEtPAIfrG79eicJI2g5Ekrctk8qmK3RRPOmUQYy
AXfrrxOVDRnHN46YnF/csel8PawkUIJ0TYunzEcBpTdb+TvlRnRUQiFl1ptfzfGIrFZHzATtfo0K
Ew1XCwpi/E11lxqGXm2VgqFIy8q1/u11bcJ0oIZtPI6Yon57nLLuw3NCpc3ARZf+8y3NhmBHtERb
p9e8qfrb2jqp/df5blaiTGe0ySqZaZ4xK7Y7zZNQYZnk2p0h4y0NXNB6YB2ThaeZfIqyO2tExHat
tW97hP5N3+qztlrcIQTOtwFnyyzrswonPR9f3IHNbROmgIHh/NUfVtZcev1KvKOZomPmAv4o3ZdI
Zg8sla7Q+Y8lLjx5AgFx41Px4s23RJAgbJtye5uoWe6BmKB0GzuJp7fCpmghc+G3SuTGbWdG6V2i
XA8QSJY16RHeqXOM0kagtphGc72HMp+ICPcu/DF3vN+63+9bO2iLf++2yXEqAJAiEIe6iEsWKI8V
8zf5MjPWB67RfE4gsB+Eb+x56eelrXssGTJ79ApVyNOzESFGCeuYtLA81pPdp8slyiIYDIk9+c+n
t644MNeAFx+OChb8Dw0CdF3eWOSjxnXgXDlX7geGiBcaJ016EmNhSMPjgw9MLhZsEdEf9GRjRirK
pBdQ2evzkJac28vFFCfpdPicvBS97v0DhU3i4pVxwC9XbcAZn4X/ZmqDjm8kWKaDIz9I5B/2uVOw
f9jePTUncycbKex+6OUon/RV7bChI1XYGv1quAHYjkzjvrgSasiDR0u/f3Ta/JnIal1z94kUlMg/
Sa6eUwFgP4srB/Ww8+J/keMAfaXR5XQLCvcK+Z2P3zKoC11gtpjrMXSn3exCaBpjp6/ri0DVaoEy
HN8jJfvjkhnN6m4jDW+cRXgJZ5R+Lz6lyVgk1utfaRU3OgUG85cVz3lI3fAfwJTaSIr2fwl2lqGZ
dxb08rY8dICdlIqmn7HcDnn4IUAsgOqSLdzfRC9kYGOPUYgKL48cNlgGHcSdVynLcoqzQv/fK/s3
SaLR7LtwPQBpRE0TRGTlrwQXd2kSYOsiMGtXdtJBWkDYARAl4w1HxlJildVjEpoKrDtaV4qR5viR
nGOh7Anij0ncOcwJei0Z5PJ3oVMGrKHUDAIexLIWlVNekmJduStVwYnjK8ffVoHM3V5djspsK5LZ
/DSSeAe/j+OHoU8EMUTY2dNkIjLZZbiRzTAFbkLMLXICFyeMtCjaoC4IpkppN8ij+3GZtFIA0HjK
jLiwwTAxbM6wGD9aqN2LP7pz6GcANBRY1/DGMRbAxyn4jZHNjWs08KgWRYnAtIsz89voHTFXl5Ba
gR6wKf1vksoDbTy1VCEsgrXq00U7Zm94F5oMDb0ou5+8kT3za3JUMNYkWgJYCyl2k75i/PIBpPm8
IZYyAtq24phNy5+RXZOJsYJlbK54tUtFdOPbLu2lXgon3ExPnh44vuK7p+6s5JS/dpsypPoDm/T1
CtlzbRxsGrCktoczpqcq1TwKTUfKVISZ0et4O+w3WtHLy32ZMq5WP74ZnIg5d+9EAX2J5y953LxU
b2cTvMlmrYkcDoUVdR1jFRhiw2knFdlslDJiUWXQmOYijxtpySbpXmm6RS7brvbgC2CKXAuFIRGD
Jq2sDWcZQOtpYLZi2YVZUZemW7teb2YTQPVXAG3F4uCZ66kWlXf3B0mlJ+WOpkx4d7+JXLSU1iC6
ZQvPuYoYaXpbBvA/+CZkXXMJcJg1EInyGUX+4N6OiVQRdhEZ9QRR9PeCP6BpIBK6zqD9MFocM7Vw
c+6QDz8iPvjy+0kW1yl9IsZUFjlGrLXlRaqb0sPBN/7k49BJ5d7/aXaXtXpPSLIV+28YIe/Kt1Jd
KhcKr93mHG+j5+k3NQZ9n8kCHQJQ5Dz8FsSPiKgqKQcibqjAsljSEjTmjCpSgEYxALAxNHgDVzj1
uwhAddJdfjxWxtnhAKYfA2HFiBgdNn8KMKsXba2ONlH39p9kcG/0IyRCbX4MP3aX6xjzWxYsGu0D
iBa6aHSvySriacRMR/3g1N+gzLvJdy5sl0q8l9ILCploOKmD74CGl7RMtjOr2gaYVhUJPF0opyw3
JQoINtBchmpobhr8AlKldpW5ir4x4vQ1rDFYswdcewtysiyjOH1yFKpTq6oJljjcCB6D/U2Tsjf1
PSrl+3+ctGOXy7xIstpNSv0zRkXwyZBb94yNQl+2VITfeNWBcPNwvjvtttp5nPGiI1NFFO/buA10
EG/3ABTIL08LukGkEEBl5CU+g6IQeguCiCByeTaRI1KpO0EMB2CPtV9pP0VpBxPgaKJz/uSkune6
Gvrjs1aXfkYAIRyKqzO3uJxsQI3cLPnasdBJde/g11cy8C81sAaYVR3dJtOhz3iqLWO/Be6D+ezR
5I58IWN8lEXX2OhT/LMC7ddKEjH0Ynxa7pvxOd+C3kVm2EQl9oLLXTgd3Nrcydor87OmuROyikhA
ppahu+LdE0f9vzTCJsSECP6KnCnnydVypj/SPQa6aEfcErFGj3lF8EreiIdn5HurKL8LbMy+2O9D
Rt7Nrn70UHfCwrEZVSB07BSTyqtNJHcsnJSvr/SCh7zuE5Fdg4yLKRFlWEGDw+stZT4lXJUfwmhZ
GAAfzDuApleJGS2/2P/gdX5BxpCdhKN+Qj7ZnkcO0lg3xTQcF0ZhTCFAbNegQUIbOe3NIss6iLKz
ZzpjPhTaElKhny5dRVM8YBMkGoM+1VBQbNp87Yr1j6AvgsEq0YlUkeWrWgV/dvYoPQLnO5Ejrw7q
Uo1gLaf2yThTaY9nurmURPQpYI6p6405vOFWoCk6nI7BFgZiUw3X/mDcq+0ZFBJRhzJu8lzS5+ub
7jCtiN84pYGuC9h5RoaMz1Qn92s51V3Pv8vPnHcjm0tz5uaoNMLO0PTclmL/mWgxI72Fz2A+9/tK
GW/V5zeB1p4R96JT0ptOvGLzxJ6xPRHLRWoSqmMZvkTY3u+XQS3JnOIcMR+RH5wqHrhsR3lVlfLi
OE9qICNzV68iHQY2ow+PpCuIMww0w0whGQMpSHyeAKliA9rV8y6E9DOPHfekVvj5dhcqwLz1sUdD
c8bQttVIoRa0StSV5G1qlB+BjPolalKzQVrf9lM5uJ2k8Kl5d95ua9zOSW0/LPbKJTrUWCO70iLe
3wlfaEohdhYEfo5ywXDI5E4PpM7FAKeQDwbYCiXRZydvRZkBw05I6qcw9xwcY/6HPBPpNQHr6Lwk
ycquFA8hDcj/EQQFJYnLtP/uXbwZHuEY8H9MW5GGRYj9qyyh9yk/VvpLeiPiz3XHBeTdcybdREdp
nTMorsEhNBh4dR8OPnXUuWME3tHQ0Pm5Z/kApqibjfZdbOmoyGb6EyX8xdqzC79/UipN79HOA654
/ywxZ0Zgg8Xa6OFUdd9Y3C/Hm1+JakGPzkni/bgnBekVjfU9n2W/78dLpzgo63lE521+UmWUwbbF
hkOEo5583lqE/Qsug3wwqlSX/0Ya1ecQ8UFnHU7iODgegqwPt2K/OrrTwQo3NY55bYWe2IcDmGom
GE8XYsnvKcvYnyeSBSV6eFHHoKaqAjuJZc6VGooL3fQwW6ZqzyWYF3rGSXpTVFNeZ+YJKhcY7hEe
d9AvLE8hEMQwSiGIGpr6s0ozSXAwx3jF1CPBUo8IVz3rSvjEC+WvwAHZY2bhpfSVrpiacH6mcCfL
yJHQs8RxaaFe008BR/FzIMNPywOd4ybCrEyU49ci1BsjLuPiwtE2b6VxoBijGxAd0E79OYujt3Lk
NLWbtzi7KXQXsl4Fc5QTG7aVPyLtPiPFVDRydbffG7DG+KssWYR9Fujbshbq4JaFtxUHzE3k8deF
PGpvMseId/CrmOJkrZp7YJ8wmZoWOoaIMjvjVPXLYzYM3bP7J98EBtGLF2nPDooI2DmPyGNFWtWq
I0s0A/lw1cyJeqJhZM78bGqYqbNSyWFWpm7ft0I6s+SizxwVVh1s/JrPLfXm53KDdZQ+jVvdD0No
Ex3ilkiKNMUkt6H2uoeeM0NYJkz8lgzmxZ4ZkWNEmX/mU6Jb8ub0IcoZFEDXWswp8VO3Qol0IGAW
DUC16+iMrY57jKkoeMeQhyGyTMb3kNq35JxeQCXvC9nm4dRNFB4hbn5M52tbM/gZ9g1dhrHYEZHJ
rBNr7MbQvYIOK0sFWgpbVUZg5cKzWuJ8Z09+nfmH4QbQWL6gTeVxsYoAJpH6ww6Dr4Zd0/zVlRQT
5b1i6HOUr6RI1v/MovzXDSVe1qLwQ+DsWu/dsHh7vM4FE1GqdBcdDmCt5jpgjtYzYtW4/BIfTAcJ
trysQ/7afCGofQAYQuVQNDrZoZxb3ylGus5n6IiQAR91S2oWqQDC6PtW8JhXHIVCt8Oo3gq3YxKZ
oupMam6s3h5fTuhmgSdbhfcQ8LPvNnQ78b8NGZH0Q8t/Q2XvE34pS6ye/R3MyTkCa6XCA8qY8piF
e+0oGn2jv/2M/QVy3yt5ZcDly7gLPEq2GSJV9eTwHjgRJN7XJyloGwBcjekTAaUc7+Fhww+wxby+
K2tZope4+i1ZoHvMGC+bnP8274iqtTICsKV8Hhxne/H3STFTXlGGKHufXYoh4hUnvMR2fy4GavSd
aT5JkvsA3VHz8OdRh72eNgnQZ7lI7JSoi4/Ej+66L9vMXtv9IRKd1Ek13IcpNaGB6Tjkl4Ve2JcI
83OT5CCPozoeCSZCbWWsXvqmMW9yM55MDoGhooifRdRG7q14PsKYwAGdwk30r1MqmwrCkWErVOHz
VANb43cXb/mDeDuPms5tLIMg6XejGs+OgIj2/vu84KmX0OGyTwZiROWMIK4kC4Yz9i+nfPXqFlh8
PZVxI970aMXOpmUHGzvzgwzPUpiqLW1HQkXSybnkrfJHSddlaYPOPT+GKsOw5c2l+qM+Go7TjV5E
1NBzygU0nA+iQNyUktnReHJsimEwq33m6cdJjzrdcnQfWmJeLMSBfMQbKn/416KIE28ssEGrFwei
P/+8wDWId0FpXC/75f2vAyGqWKdZ38WaQ1Cyw3vf15Shp2Ng+n5gZpkUp9LjWCcg/qH54Vu7a6I/
3D7uq+v1LBhLBwN+mGhUNaruFN/oKpKPtf45N+HRDv/VI/sS9iLbFOzEiUuYneWlhJm5ORGY37kj
aszHfKdGYzV/DyqxhincXg00iS3pHzWLES3ZZ3bVSPSkQpKpFpg7WBSLMJWGfH8dn6AcOM+RrHsh
GnLkRlkzJ15J0tDM0keXT8C2wAEMQXv+1l9EWy+xh3I/FamPROwg6aAiCAAplGnCuzT2dwtd+Poj
3jDSdwVZ45qmQgQY6cfmOBTkxHU11ivRZ2hbJMmM4PfstnkqsdCIOqTDnLgjzejJVz5ZEh4bRKs7
I0IG5odfYlhay6pymB2G3CQu0ejeTID9szWNEILyPd8WHQHLOKZ1nsmejUdS6eLMpDyywhfI4ljk
mr7NvW7NWs4pcKQZCGk5X3vLVW61GeBfkTbyJxfvIuixc/W0LDTLJjSsvaGm6ycu0oh9HJ+75q5y
c+ct9UtgSI3NqcU3Ss4KD61d+htQlkhZZODjtNwBe30agcM1QHpjWn6LjknLIXVyxRXkeIjkpWY0
KnGMUEcIK/TjPKb17KLmnPZ/HDBZEqpLuicVxighGKVLZaZkpuqYmxTEg0uk6Xskd9+aMoLb2QZX
GXS1IL5C69EnbF05V5XmsJhFkTSo543PZqn2MmLdyDaEq5+GNx3cRy1LwbFUFniDKeH39DUMPZOe
PtsRUjFc/cG5+QhGFgp4e3+JEwFvou7K/V+AzLZiAUGFecXE7tVsB51L0O7SKU4Ik/9OGxE+0Nqv
wvQy9DIiQ5B2j403W6wR+9cVhliaiJf18fnIYU8fUQhyIOheYoMc4XylOyaHc+TO/yGeYilPnkMa
fSJKSPkvk+tTaWdud7KPuh2xGvjv3dncrtBmDfaWaXmum5tb1XKlrh4glOQ/vusr5jsaeVff+Lfp
IAySAw8cL9pNh5O41FzM62tjiNVlIh5A4nb7YS6Jnb05H7VxPlAuGhNHWV+03dclne4NIuT5Kc6T
JbBeralZi9Cc1kGzp1YdZHzMjMjhP+ozfCnP24T0JvL0Fvp1ADSPxU/eCICNnl47rPFAEO/LYoxc
hpQ8COhjPa7IvjIZs/lFTgTLFu19V6U62LEqK1j2NuTuMWCe38dApmlupGRpLcm7sIEb/3kL+Pr7
S5oU1xx0IluFI89kydW0SZ4nXtQtHQxl9REwvl0zFawMrsuZzK/VDpMEjXNTiSpl3GDW2AK4eoAk
aXjOrFxzlr3ng5LQ8uFYMEDjlQPxb5EP6b4/ZxZHeWD9pOajVu9c16j59RPb/N/Bw2o9Bw68Y87l
7INBq/6ezESQUY1wGOryQgaeDMoGZtHJgp2s4bC+DcT82LXQpT8s2tY+8i1XDdO6X8REfrNy8gCx
3VdETu2/c5/3YGCGxGH5b4FeM0hxSS72plOT3MGPNvXKLHmXUka9y6lyIVxOvZP2WkM4ce1Y+3Ee
pbH5F/vjqKW2pEWRQvyfQ7Nlgp/EOqUFaL2zgiaRKnyTq5Y32a0WyzkYvFgdUqvb4etH5KMKzsTt
wpQsaqnMIOpV1IcmK7moqH9bICpU9LFf26QwRgFFpNtFa7ryTGi5h9iOOsT/NhENbYtKOw3ivSW9
POkb9lAsfBxuva4PJ/jvKgUdFtSTeLvnlaERjBnqkXQOG+oGYb1xkpsTvW9Pce5SNiffnmHI/Biq
HF8Kh4ixybwq35RBgnTqIqV8YaGOsXAbkbd7fktbywIwyZQ1buthDevfxWWIcz2nr/vxA1bjJI3m
sIxZyq1SnnTnbLUrERDq3k8/d9mfNF4vLFPZX0V0M6w/yR8pXth/5opxJi4yAqmjoHyNjVfBKWuU
H/k53/+6IOETnoYXE+gHHnFjgWNV7Yv/HLp82pNc1kLShS+pQNynsZbSR4ULKgad6qMeD2a/isl1
v0Ns73Lvkwa6Qa2NjQCiibq64OUlbOzKfpQDF2vDirlXZdspyQEcIkp9UFIKKJZEF/Ig6NS9zwKn
BLhr/MtXSNseKPAC1fYzc+c5OheQzQQCmOOukvpuwWwMdnMxtqy5DrSjJ0CbzNyH6j5b9CnMhsnS
icHGKKqlp1MNEObG8edpr/W5o4PqUSnSC1X3EEWSgFQPdesDjciOmEPObjl1ebyP+E+L2gil9e0n
OhHAcMnWDX5p7N81KyUuyy+R9zHfEGlbuaWqtAFUsefMxejYu4Ahcytwn+xIbQJSTIDL54IOcPVv
tSpENubOYNx1zEJ9QQVnkfifiv+5jv68crztVrbIfhQo4PAZqTWBmxxP7fEJSrvjr5ffHT/5CVE2
r5+LJTogkKYg6atZzBE5KPWUsTINCILPdT9ZxICloW2KJ6pBdjGd9rAhPS6j8S7Xw6FNbf2uuJ1Z
TItUjGbWOmx9cQDDwGN9m5zGPRVrYp17BUjzdWLa4GEpC65FdM3RiRuDTq32lOZ9RcD6RP0X6noE
WgMTNURn9/FYL/Ke37XaebdWQzfR+eewJlK0tSyyobjpH03x6UKlvOs98AeaFhpWiQQGZgoVo+39
n3vShjTMBvaYOBZRrsQV3v4213NLVjT9h2fYKM17Nr/TEli1bNJ6CTf22sQPxTiNffVrKC/8vHuu
x5B/B8ZwjYnyHEHemCwdj8Txtu9eG8Jib8sOBaGbHpg2JQQUAMWHJrdvInZJvqMXEJd8S/wkXy+0
hzYJ/j4t7gazdMd+a3mPvHIMZ50xIK61DVhJZMzkzNJpjfq5IXCCLlaIlHkAbJbnbRVcAYUGOddW
6tl/4MUUs79vtiKiCdcYf4gMKsTVHQEK2rIbVcu6en91XfFljMtqGjYzj5Aa8D0gUmyAi/P2O2eW
USubVL4WBc8egOgqhaXtepxAoCdiFYeAetvjo41SRscKzXJI0u9O/eePLjLx4Fh06Oo2PYGGwYxM
XxRrKgO9A4FG7SbpJXA2jdEcEG8MFiI1GFLv0guEKeq8QHcxYwHewwR05pSkh7oi/03m/xov2KoP
+OWefvf55F2FKCWi6Xg+UFg6JIdaEq54r8bTLLm7sV8AM2oVj6HwadOxpcy+sm7vSv0gN4Wh3OcX
MPHREP0Ih9OOQUAPZwZq93AZvHDuk2Q6wRa7mVOhFR9nye+011+6Wr5ueGNOnQ3I6j9gDMp/wgMR
DCI5RGFQhJCiJyRC1Bgq7Vvr0CDVDsOYhxkO50pRg7N+qTDANMxyGb/m3TzxAR3ghAMhz2Mlib56
crFpp2OqQ69B3vjjFGSBbCR6+maFH0U8apy7M2Crc4O7t2ycnlL4hY2VoxrRoUVxjevEPIWGU0QW
sSUUKjX8WHvGBkCWJlxvyGmJvA5Cnq60hCBlHoUKCUi7JC0T4dW9qy4RrwLDKvCAcb4Xt9+7H5LQ
zC8zfF9TmV0JhNeY5SmrNsAV4ZqVA9Io8qZY9mjTxjMFeYAzHl6F19ZRZleTPIrfgiU19K/LdQE/
zdKAjsI406Ue2aQz/Al+QaJZoRQAcbfDddjfHIpwSve2MQO9q4tY+wpbwDx1FlPBfjxozaa3Cidi
xkP4kdAPrXrDrNZhmYrQj6B3RFrKne72+vqaVzrFwMZmD6LdKGF6/12jpYa30Bwt6Zno77vawi+s
l31eXHwnZT++3nzz4GAI6/cILKSxkZIfiUvv3u+UZeAuLCNpAyne9M05hxMfUw3l7FS2V9NATDBp
rg1ELnGO+bZCw4DLIIGCGkhJtdt6gEq+pkUNI+j+MFvV5TG368WDjdOcDri9WqlOSgjSuP4rIf3C
+aGyfDDtIE0Ya2HoxKIlBjzsFmEFa3oUlD1+EpAoWjIuX7GE662nHaO7xtV0Jdf9+QmCMTUQALO7
4hCZRgY17TCs9/HtCIbgqv9MnePbI+HaG4Sj7n2EIEFYGHi746VlRqn5N0KX9aYiy46FoHfWhhlY
4l/gtjx/NHZMqkRfTtpNlEAH+60Vgyv+CQoVdAvoHVCKCeXdgkcZDs2Z90pm79HrABa9k3lV8sZK
xxO9YrqUbv+sV5Pe0l+c/fr+Bx+YG/yUc5E3DuPzVBjErAa+3T77eUultzXC8akBi0nnjq7zsapK
gChUO3EteP9yFSKTgymF/CAppS+t/5EkjSDsw9k0MWV1k0RTxxl466LaY00SUV4qf87xJAltBL/p
zatK1jO25ChK4oZN7s0Qedlzv9yCEBGQ9JEIf3RJkDPIszchaX8CX7Am9f3LKVM+ONziwi874jgG
0HYR4ELrqxbv67OEvUnln9W4q+vf06Ie0BoNrKFktdGi5ztnpGLoXI/xiAKI7cWsKoCyhe9pa8UE
jRpSB4QrkeeDzrvNsnwzrOoC/0Bc5Oofe7YWDAoB6AY8Sh38+xfPH83XhrqMeTlje1LvsJgR+OXO
jUc0ra5kU2Q+iVEh6KOF7LiKHWKOGavvwpX7TcVyLdBjVnIfQVIOfiISIYs1UJxR0rbfNccAW/gJ
fNf1GI1jxzxvpRO1qPkKcWYs/E1DHw6XRqYplJb65hSuZ6mgdOJsCA4+m9XdBoXb0G4ZTc/IqYXx
BLSwbLG2/e5quvlEy7zzoivyLRN6fAEqz0tp2ZTg5UUZ1GJ+5WfAUBicX+vgGJiVs0TqInxueeDg
MxL9wF/Z5u0m3UEBFv/ab0ZDsxmCsz7h62ar9XM09Bvp72M4mdhOzpXw7D70Rn4c4kLkpa1o1/Rs
ZUUdZu/M2Jog9ENrLv2yGYhWvn7KzdbfasW8IqXzU/1xD10IM/YqcLUGby7+DAKrwkOmMoEuL+Sh
/GHN+lGp9mcxtx/Ea57PaRHaTATyFBwsCgNt9/oO6KonQjHfT4A+ggKRP82C79Z9WHH7XNEhprAn
kcuRgLtXAUnRM1qRUeS9EmbSMPcx1oDAq6nbf3l48QEY9nMnj15HWI2Y2tyPIftZCxsiHjK25Gu/
ibttWbZapbIPp33Sr2AHyyc3sW+aW04j4orS/xbatwYObRdTLEjJ92kwjWts7m9Fz/Abu5zmngor
suk4nKN0/3aNAQAKeMB9YB6iZWzQpMe28cB0AfmB8BPgdOlCz6iwBYdtR+vTghEwRzFSru4hles9
qzYRuraTvDi7mnYOEb4AV1osO1z5YsRdBLRUMQQAkQYGYnvUTONDSHgXc/Dtu0O/atnVX2CXShjO
CW+JSpDN4nYlmF5aLNsYWlK8LscxtWc1G23JjByVu/DPFZaHaAJoi1t/4XuVpxByUj7KOebc3F+x
2WWiig5X4jMQqm+nsIB86T1W01l5va8JI2nCmlJFvFRPDh7waNAvcAmCrDknkHE0ENf/5N3tI71a
IPxs2fOWk6B8iMk8gDmfIklpIdP14tJfIQfdUto8iqLd/ZpT12oorPvvVyni/2EvNRiHUMPvyzDP
sA0BGcZEHdkQX01w+io6vNSvsAc7iv3Fyic5VzsYzdRyoFDengx0BNmWIuzcagCzOrhL1oUkbz6w
TUjABExZVPuE6Vdp1DCrTpLDDWLzEO7q5uxPHzMIiCgoJ8sNWY4XMYQcsXZ9An95c88gpdnTK1XT
aq+2gfNyRPYAnul6tjgpWr2D2wQ7v0N8rUmIzi1N4TaHrTyP3iMMfgdG8dDE1hd4k83+NE4RPhoa
Icw/HaqsePuMHtaS1B8C86Ol5vfwrFQUi3168NfM7FyMe2FQJa1I17b0vxqoUAU/OjYhD50bVoYJ
BTk90rD/L8xOh8P2VbduZ8EvFQylm9zpnrhFvlqa4U2ssYdMkpgRgtueEjbqJZSzce+tnGEAuVxK
luXp8oRck0Rt1266wkjJpeoiZmJOLvHoOaWjSAj7f5jLRjs+pO5CpMS/zAPIJjvCISSDc7ZwBMNR
wBfSdsoqH/Dh7FjE8cy94LUdBBwp7j68F7AavxxHcchJLZz9MuHSU+OjjAHozW32cRHSPMPIcznu
8txHaNmxd8LXwKiqGdaK02C2Vd33o+eKp7/kJ6HRGfVtdOaiVlN3bDd9a00/rlXJ0HFartZnltQB
Tyw9r4fbD1VRWQkFRzb/yexED230JM5oiZIMFDqwufMSTw56DNc4JB+KPwRK6XZXRgZuzXVSiXcc
Afo19Ktd23wAHSUgw0zZZLDs2P3W2N6oPw7YDnELa6SNmMNmRzXxPJOz32NSbdKvpbIt40xgFqaK
MX1I++zVdjVWlXwdcoSxdcPCQNmZWIIdG0ZMjBjGyfLPNKgoG6yWhvv+j3a+FEANJ3jRSGyXTXug
3ID7CySLmDqJ+iA2R4KFcS/yU5g2pdBmdxlX9gGb5gXFR+wzFc8xDu5ng5inY12O2lhqwryh5P9o
3mm91S4386evjTgZmSOJgDUd1tv/ikY5i8LN0+L5+ZJGLhHVGDDX4kjerzgyR6+c4Do2bR08JHv0
fYFyTKotGibP231pfjhUUSP8gN77OXogIEWsfXp5AFUJzoACnlq3LqwOtkJRpYzbtypOxovZ8W1C
1nKk4J3o6wFDKCcjFvHie8GgCGeMujP98RJ4BzipYGC0M5toMGR5EoOYACDMOUi7mec8mGcZo9JD
BiPiV4YhItk0qSXWbLskVevBuW+GBPNlknv1KVCVdzqQmHQgxiWgwlJVi7dMlBjBzh78CFfaHYQN
0rC7h7RgxvOM0HB3mGXtzD+NOzv4NTy59zjB+1m6JgRfKqZudZf9iBda1a1dU40006rLzEsJ5bgn
xm9ybBrUnvtkgEmklXkRZlNzXggSitSI+Y1sm+jq3SZ17zxXuazdTKz3nE9FwMABl+dogTwxy+2O
cDYztSQnokfl/s4Vsv+H7VPgcMG5N1bZQl3P4aLeS00A6yoVXZ5cUBjCFxFLZEXFqQvlqjVpbE70
dL3wU9DdyyG7TQcD1ZBrl8o/cyK8sxtOw45oeCvmWQjdqOe96voOltG14wS/hHz2XAgP5YlgeKFG
g0VdyMXy6dCLRKJFzVKjV9sI0NYiaacMO30BJrW/ERNtDhki7+Jv2T4z9aTNmuVG/8o62J90G84k
QGYFuk1bGRqjzK13UsxiiV4q+aWiLW3j/Q0iyVRZUquALKjNILQqdRzSpjC/m0APymk8BU+ks26b
6AQ5bAtrTviHfX3xA/78BaX5dgwVshR08jtsjqxpKJ05bHdoKAcHrCtpl9mDy6jyymcIh0zIR+S5
zyJiLCzd+EOqbj8lmB2Cg7BmiJHO3tXUcjDhzaiQpJozcUJnERc93evtkZAUkXZ0ze3ttPxTdk5u
CMikGTR6N7Rz2mto6cYTmpCiz/Tuo7OTVIGnLxTeIzXfts+Fl7PzyoN91NyM+QkqopPiqrDgo45N
BuUh+0bm2M0HMHnnh2FOObDZNz6Uh4I+ntHC3Ri1cdPPSsljCL6oO6J7wfMRhGg1CGxir2iEqJFC
Rl/5IE1KS0TEHCgq6ea7b5RwZCDpZdqP6DN32pdjnu3BWoa85tyPn6AO65AAPJAWbGb/s4KkOBLJ
ftHbl8kxWG7/46uui9FhYWHspWTvmueH69cyQ7wV3nFlZGqXL47S/zlEn3jyaGDLKH7fq1HZ2T0Z
TpGh5ea+cDj+xxi/E02lRcCJrncdEKp3awJDkhylQIpsB1ASsVBZfZ2bfQvmtTJS6SMcvdKnuWQ0
ytMLr/2k4wByCwec5ZcSOHlp4Mr59OYgHXfOvkMdLoc7f++AxnbJL17p0sUyojepJnXhWaXjeQ1f
ijkhFrTClFN7nGtrHkdB9pP8iLDFtswbRxGAu8ZUrkuLPM63nrHHSQ5kXk+nGnRyzJyt6m27fhGa
YA3mYqp3aRymkPDRACMpCKlJZjeSLQxX4lsuct0fdNu/CXotnsfZMY5ZRJJAx8yIuPebUA0jAecN
w64eGHOyBP7j0zTgC89G8R7967XWcwRygCCmaUb+oWzujIggqlzFwi7CdrjdhrpqgM4jFdrUzxp8
pO4kqWovFWIVTsdCJOVb77TDXnq+5xgEiTxUBXlxQVJfuQtrb/NTgha9NKeoCRtWhEL7FQI6+9Z+
83/pIsorqFU5zsDtamS6ZmScQLyAXcktwtWa/RsUmnmzGOsWfYWa7hJCryXvxyQ7VZF9W7yepGzc
UvWg76slKbELDNF4hWSg7ZJQDHS93Z7TflqHUqXvw6VVoYtRsniJZaCDbQVdrEp33PEkGpL7OoUx
ue5TEE/Nkilnq1UnQqQC4XVWot1cHVKe4N/HiHIWTp3IG1KlTDLrJ3FQygVPt23Y1XBlnhLWWXzN
TVN30N85Bsvp25M0HTtYLQagcl2LVONwd9Bgxzu+BF9tXTeLIhcXq8ZrLft5Z4XSug7kwDJsaj1q
vP7sudoxlBpvNQ9BRpoz0rdrvW8OFYWlktg7I/VRm4mYQp3sKpJwxpP2kgky7I2yyH/YTEixe+Xw
8HiH8M8E+w7mUOVvg9L7MjFv9suBPKPyM1t0JtwWtN2ocKMcdqt6K73RyZDE7WWyacm2ZX62G7dC
9xpSSArzx9qqhqU1IgYcEgqTqep/YRHhICqgnVglFsKUFbPnsQqQqM3I5+4W4ysKFCwMIt5YaExI
uBrPx/nVlwY3iRrX5sfdfywWCvHpF7ShvvzDlgMA934JCrVnUz2yQwg+xC8CjqEB+VOuvxJFiYd/
ufMEJfBJ1D75DyAySOQyYIIjIj8V1o1NtcsHQj50i8NLPN5KwYF+YEe+to2t3pxTt7wuGRoFGOc7
LdmCMv8REsa+TjondFNQHrwOMaX2k1enllTUsiYQeDuxKMbb9L1dosWsCNGXVcL58JCz91yYYyoG
w3VE2ao9dKXFiB4WlHFJCSrHk3YlgpL8NL0urZqBb2hlv1boTbOPbzE5ix2diwQkBsDtz3ValEH9
4RyGMdu9xmF18Jt+/5ajlA2y2On3pHaUb6JKtoVBKk2qK9PHkD8c1B+7CLpQgEgFTjDVfrHvcuSM
6A6t9a1ewzLpp42fcp9cfz5ilAPajLlwRE8yMhf+b3FddN3RX7a3dyYfk/M5zUmNgJfkpMyJuDq2
Jx9i3agsNOjC+Zb4qdazOO9ckmMo3WNK2GeLzUd/ZcicIZVSD5EfZ5fXnM+2wqgAJhFKamYFPK44
PoZb3jDtIH7LJBCaUg1A3nt/lw2zbYZf4klVM/yS9DuJKCkNOKRG0kDHd10oet++bi9eRDA+j8hv
DOWBSU77NyR5J2j2533C60F9T/nns6QtRHdTAC9BCU08hdYOGjtlkcevscwxyVNxDXEwtu3SB3f4
+peSYQEL8D9PxhjuYXhZ12g8WwgZ/iFyuP7MybfgBKldaYbM3Sp9HExVdht0VmTh12j2ibQpWxMy
dbTzJi9Q2GiXR4wdCVPoathX7yzu1DcIMIM4kFEg3atTqrUWVEy/OQenyM5CFWJSF+WOyI6goLYR
rHFmteAjN6J0z7QtLcvYpDVXUwOuTp9Nxlm0SODH+TqNZUDh7OQ7pV86vNVlccKYcQuIlkx6ZVHw
wMMoGcrWUOuMpm9TfJdmelUX19ZAClx+l9uwEl4I5eqFvkPgq2YB8ogg3RZo0vhc420PtkJMxTEA
fihOrGDI5d0b/pYZu0zcK8yP8d86dgkSPDylapmaJpEQz9z457ZlwyGZtdMfrMw0Pw+a+cl77gon
/2c47driBq1NmNZJEZDFCu18KtHpelVkxQvGzEpCM/TFJoYNBajxiFS11P36jeEbLrlygDoeXIN3
+2IbXERUlkXO0nOPRXJw0pt4z1XS/WpDH8+1c7lKuIpHl10f25+CclFDoJufgbJNKFjJxuqElmq9
3UVoK58qeRb5CHbZiyp2h2hZtQfUYO1l13oKQZ7G1KmI5h3zKPGjHevxbvlzWGYHQ+wEf12GGcG0
nz5CWJnQ4SFtM7T0Q/HQldt/WqkAeov1erlT2mNyN4jSuTHrE1shWzB5mxc0WmqMewyQMD3skG2t
pOPwhzEQODKVW42QaTwWeFKD3KBFlPkOP6uCIGA+FIHL1RCp2LQljwZd/OefqTeYyVIKl8a6BlPJ
gUsjsFevWHitzkRPhBAtj0NYgvfKBbUs9rn2hqlqe3xhUPUAxTVI8plZsYGqkP4+3wo2HWAX7aZi
dQMBKAzK0zqSPDCuA2ZxVzGMO+NFlJlZ2W81LDhAuMvtnzSyrUeIyaduppTKRemGuDrQ80W4sfUZ
F80oscXsX0sJ5xPBwYGMsDVV2EHSlZwqvMBB03ZmnLBvCr0pDGTWDE8DZiNx/AJCNdVHoB6cQhMG
/e/jQ/YPRNJrjfgpsugSp8MtYQzVigKIOzA3x+er9754a4eG4QFA99O2SaJNRg3ltrm+Trwy5CMT
9KifuTKO0Bnn5gzE3p+VJ0iEQd79rRbGZSo2RJgY+Y4rOtZ1RKDgcbxU6gIMOHzbuAqBu1MUIh4n
8Z6KjOrn173DdVSCOU9Tc4wHALW2B6rL6fp8TQHgfvcLJHA5YBry0nU5+ZzppDiiWLrWm1phKYDL
ZanJ/pEyPyirGvr+HuBJYc+iakB+IcJ1ze9BqZ0VpfbV16fH5BOJ90JvsTBucZxCteDKk9C5Pj6j
rcpBqfuDcdU8iCmxSkBPNU4XkKqLqtKEklxfiBVT8UiOgKMM8JlnCiGNI1Mp03Kt43Mn/d3+Kt9U
83cu+siKcXQF3BhNqkUz3AM0BBMGsmJALndvAH2Kh5/5fbxqsn03J4otqf7bqE+cjISZwh/Whm/J
hViqaRpVfn0iaQLo0RwHBRBNq/dcmg8qQLCrHOT/JFhu1593yEKnAL9oKmGWBoTQICwCe7Q2CV4h
wJxiymUz0voyzRtuoDNMAE/NEoY0sajVRAJ+AcU35jRbz9eqJCxRWsofSn43IvFAzyY5tIqFBMux
XhDyrJVm6eMQIvpasmS3/6Cl0qDRhJXXBDEkao+GSnPpFDK1GuJjxDUGDXKxDtdr3i3PR/tDNZ9P
nOw5/ULtVoS9vHqram19+1oWM74yvCZ/CxC3Ht0+z1SBXY+OdxOyan8GvY093BgLLUfmfc41JY00
w0UWQ3qqBomn24Swdw9cMDdJLXaRBPZqnww5r0iCBU7ZGzWfQAmYPXYaLrdoaW8y7d8WxD1ZiYMS
1AVymW3XYroY1yJyl58vBTcTTtM2EXiKPUeSi6I2Cg+zFA21igD2jlJngkezV82XEMJU0pUx8iX3
MUBl+jrmGhvmEMEEWVOZeRYD6Aelnn0egR2kgTzcp2AtucEMjCdorn1wUQD9cCBY+if/hylFTdMz
7PgXNbWNoTmN4hNd51ZPDx6CgIVwaAXI7v0cnzKGUgRS398KsU3/UdjLtgJSNtF/jwviRHCT+RB6
QV0wyAgO8ZyIY1nlzTqu0PLww5peDa3xk1OHqPFzs9UKrUgT+fLalSV925KkpqmUsw7Qxn3rpKF3
5ll75n9AcmcGiHsJATuZiXLhn9rNy9OROsgCQiAKGV89NmbiHyVVOQ2qHMFBMB/uGMnUjo2C4UXb
E8mPWP9IBfMZnFdqRcM/qiLBHI/RT+5YYFI7cOt97pu32flcwDnmlhK85bgEzCE1NauGlkPyO6Zb
R5fw0D3aOMSRdZwA/H4aKZizITXmuHUEGxKq9bbEvLQiWW+HPmGauZ1BMMNtlvw3SVIr+6UXMZH4
KHtXk2tRSk3rDhOSey2TC2ZpaBIM4PpcyrJVu58idqA3ribC0xy1e6URqrPT4EBC/IgQgrFP6+TW
NgKrwSfbIzq0xcfKNDTsE9ZeHxWhTUzgy+LTg5qZJIjj0OCy04DnjEI1CibcRyOUS2q/fkNHJ/vn
3kVTxKcY1MtgGI7mt8DGwMbm2ZBNM0YIYwpK5H0ZLmCWi61HU540RwzNCca1H0hkWBDSE5asD9aY
7+0JzZqjtJhS0zh9DLHHOV9JAem51ZMHvSM2pwfz25yr+W0wIotGdTWLPY7hrsYcjwymOdaZG2wh
z6aHZAMRI1NNQCY46n2Z6soiMVoVQ69xxo4TguRd2tGh0rawCcyqK16n3fJQGnUovJ4dCV+wU6Jf
MaLpJZa8l+Du/SgtYuWLz4snxvgy+OqhC1ki7VCmk/VyV21a4HwSzDBMzBkRzJZE2o8gd/iYebO0
Xis8MrHvkAKW5RJueXxEX2zAXZ1O6QIiTRKeJgvuL52mi3wa/LS6Jbs8E/H3PVNE0BOwQafUOKLg
0/yntZaolov6bc/Jkrt56X9etJD2V+CNn9LrJA+ICQ481K9X3KkuI92fAt2ezR2dJvbeWW9bx0Zj
WU3DYLDbZxFLE0OQShjue/lHECP1K4D5L6q4B7xFbjqdxoQ3uGpEuqpWm1Tz6dFHJvcgprjvWyAc
UAzm5nNa3vAaGn1hcnjd411bjk1R3Lxb5szb4mBw19Z5FH2FscipHeBSA02YKsvql8EbQ9lXKpH9
e/wONFbOdhzwUCOCoSlw6vn2eCdSpsVDA8lDLwOW45MfUMg2FTrCsBM/HEE3XUGyNba/SUwE3dXj
AWjg36oLR4pS3UR+I8w7IQZK5Pn3HixmwW42UXKSbnhBEpSkVZZYwG+6MAmZk6eGTYDrcb66XsZp
wpzEbroDtyWVXg64pb7FCDnVBE+schY9gXgQllSDwwAd2SgfQ6GkeyED8BdbP3JiHsgTdlpE5m/c
o4P11WjLvuykM1Mvtu8DMDxp/GUI9n63RrFOQDEatJ6ybD5Ajh/6Gx5ly6qyDpfASZRcsBY8G9wf
6iL69qefIQ/GbTG7fz7Z9Uu3+YzdfMHve/cabJGH2GU2pGiGFbaw1vzMCy8hvQy0ksTLHamJuwps
C4kp5mSKQBl8jBo3Wl5/eooZpthMY3qV4j0wWva6Z5BJ3rc51i9X5Jxg5nYLJ1qHMkBWcGdRKGlZ
RdjcIGmuRzkV70FgkYmCHrmevlP5IGW0RQSi3oE0M12qav8i8/cMqz7LlrTqZD0h8OT0+W4Buv/j
5J7rR/aIyB2D00CCmLPkEDgGkXQC9PMUaXHxpviioLR3A/RmQyDBqZs/dqqSfrzsRcXd/vuJq2jm
QFPS/D31aJMvBrmYATffo/unUSUTCy1EmZ+D4GzvhQVBzBSVerQ2yJB7t6D5dMOqMLyHJC2AganZ
rDY617mX2m3TlToaR1FgwwDf8TvBvAXaun0vc7QVk5yirqsVruuq6p5VQovxUJPQryOsKxF/ivg4
q/06ssvnH45uZYcrLlH25SsbFp355j4/xFW5m0YZzrXyEEmuwEDVE/zAnUSy+Srv5kgeCPp/kI0i
/c3TNHe4mgI4iaXhMoV9C2/gKHQtCJsDU4Zx+CR3DECUDoLm7cx3i9z+k51c65QynKAqHzmrJyuG
gZh6MqQ9Krx/dzsYCA2DnWn7pTETkPRGDGmvpp0vSoLHESFBX65yzVQb+Nge4j1KP4o1Vsq6FOlf
uOPrCeUJaf3mz0gBD4DS7YoPp68gCoi3oZtXfP7vc9Cvu4TBIk7z3eFCAk6ykmd8P7NZkQqObVLO
qe+EHb4IRl1/hRrV+EMF0kXegvqzoCeSeQNjTLMpxITzWpreLajXM5sAbk6qu4IaRJJXBPlc0Jjp
NoOFIJwrwD79lO9rxjXCwkZUBVSTskToy9+wFQy9A6+pJUi8VoMGy8mSDnRLr/bMNqmviwWK/Jfr
aYGfxsLTo6KJD1Eq9Q4q4zPyZA0FTW86bBFLEpMJ/c8zi9INGWBTdkRWmhvo2uJq4NqM8Upi7+HN
wk3wvjSrXIA3LT0dup1hlhM6KvRlo1jt7p1AqWLEGEXPAeEwgewfV+RSdII5T2A0saUVSkjAJWgP
Ez4U1V0Z511avPgOjheB1OcAMMMbqCNuDQwadLah7BWNZBu9V8n38aIPMeRDGlMTHPt10S6YUUTB
mgcN/TytkGnWrlacVsULL/plb7tAY2yhc7+OzyVvCl2cfDjXw/YQuRifZfdLjYB18s7VoxEZh9Aa
zWJfVqw0k7Ea9LAmn1D0FxvqFaNyI+94d7+QvzfBWNE83RxMeec3lyxDEa3/8DeLBOCXP5zqzVFb
vm2P1oZFoWEjk8xvwPWc+L1K7bdpHfDt9ppJymPqH+LZhYHOgVGA/+W9iKz3fRcrGJDugbCplgr+
Gcg8IcHTtgUTG7wz9s5XKyRhWDdwFDJKDQ4DjQTtJwQtChfgWFXJDvkAesh1UUtGPRQtmKv3Q/Db
6L6Jc2ezktz+evRB6GErOulanMWCHz6W6GM6Uke3ckA/2FYrlSp/jOzYlPNhnXahrS4K12cRzzLS
tybC8HPLzii0HC1sI6gbJJYb+sAMNFnb1EkO0F0nIxLX8rlD81NT1/jAdxL30rpAqroiBzoSfEU/
t7EvJUE+mOYA4UFlZYUTDNZj8rpe+/jpGaOceuW54OAvpyoCTWNktGZmi8MBQ5KTaIW9H5InePwq
GEzms+3Q+0HeE94V8yw9oNLtBXgwSwInlrCytgGdxh7caEBCNOD/icTwxEkPPikvLuWn7/fyRLPK
gnMM+s64VJYY4ZP3oJ4yaHW/s6mJ2OQ8av57phIb4IN0uvrRwI6wgaKV8QHXbxdikj0VNEWxORFG
I1GKTIBYPMfQyRjwAEJw5QfRW/Ia4WEh2qJAP4hxw9DQR/EG+SA8I6JS56opxvxEbb2FQg6XTzc3
oeg85tlk1mYVcXS/E6cb6oeWPwnuUPhOeq04TNZ4qj+Ne0uezhjtUQTugq4qJfW0dGJ8UEYEgM6b
+XP8RpCRHOkH0DLWDOXO0zUd503SQhCU34eCIbbLhIayXJtoqFdnNTZnMkK3mAWjUK/iFjfnkwkQ
QU2UTA8mIaePKICspHf/YAFbwH9Yst6emb/ATcjUqmg8ISvDznAXXkxghDja8g4FoVx1KcQcAmgC
o3az0bmgQqNgPjy50dHx2fxjNbo+M8xuCd/6pzZvzjy1JHR6QVsz4axiYnCMEf/YS4PPanf+yWfV
lRhAQ+0ZTKD82nFpQDL4gDqdKB3OlR5wf/ZMBAjSUjQLhFiI9JZQl0JRi7TT4Jerud2vPCRLdeZn
pDVHlKI6NrLTHF9dr3k8ooS2FswyMaeNZ6h1SsRpxMvQ1VxZ/0HJChvnc9s9G+i1xnwfQm2/XMbK
N1ZiMsz/09Ye5cOaHTF2YDFP+FvMKizZTu5FuVUaQcowlqsL9TKRcSqT5ExYR4ag9Kfc6ergW8f4
ZnlCGf6Sg6Ii0zIzurFlTDNKW0rY8G4ujgBzeKP1MILKpxzYH3MkjUoRBRF3KTMriEtnVY6vwCpq
Msxzsn+JGVYXmsnJiJQyBUJiAVHKiMrKvcsef8HPaXwqAQ1517e9Eglv2LX8fx3h3dUilynR7ah0
F1xwQn7OxjWgN3WRK2C37qaFTHTkTMU1/c+5PHBzB59hS4xzOGaMzMLEULJjkHKFPN8HAc7NTRjB
L0NdhHIUY5Q8ORLNfeblssiUA03cfi8F+iFBG15IhGLtC04RzwhUWCUdPCirwg+puFnK29QXTVUl
Ydpn9p2LkoIIF/h7A/qcpocPXxk5e26i+7zIzmiZAIx1b2Fs24pIk4mgbf08eznlCav5HarEWd5g
hVflAjVx8/Aa8TswmWM/vvyq6B9rD2ozodvL8HlX4s7GDbcW1BYjauIrHr0zJ8w3vbKraJ2XNktH
cwydJIaXtymz3pDUroVY/xliFFuI6fSi0x4RIIblcIctiqXyHT9MX1HifSLYnaCn12g6n2eqdBNN
+wYG4mz3LTeSLMGDgqXs5c8HycW0LzRwANcR7bsh/nGDI/3noMaUuJ2Uj1QVyHvtSMSSh+I6TVPD
S8IYWRTE8ci2hnd9e+oQUMrG+g0BGWfbmR+klKJlNoqml0G4RH8vpDQqoU+BYx6xJLvhs+UHFDS3
t6S7Fht1JZfmIUPstuzfzn8qjx5CoEFtwWvi5XT6vY+hx8SageWew1Xd1itHoCybGB2+guUIlOus
25odcan852abp3xND1nhl1SlgAnA1K54MYVuIKLflDcOXfPp1QxAqDUqOIkdVz7iR2EzAANJiune
H0aGymiYeWL6UKLf+jvvkBDdRCKBM7d68gu8J8VC5KOGriqyZq6n1iMDjCGxNXrGwQb+HxvaX35Z
izbKh/JNMf9JQIK1iQoHrKqt15u3A/NsrE7SxslWo4LTShHe+dlhrn18WEi7YyWZ+7lLIbdT86jY
vm0u9qCfdIJEXueP9OisWERiwExtexSX4sWRuAp96De4J3p8q9OjtrNdVPuWaVJlUKZZJ1DH21o6
eaI4wDNhBoEu4KH5liBETAUbdMEX69GiOwA6zKekj8J4BbByNJDYYIb8e9FmYB8J9uqLtf5DW3oQ
HDE9ERsxOBMVqbB9irqVo+f2LZmf843rDmxHeh0+rS0b2regVMtX+mDI3cXzFSLc4E3fuEFxz4/9
ODp2OvmJRR+YxgwHfsDgmnqsk2jVk38nwkPwA1/Cg8Mz4Xq75l7vkh9wl6xJQo4kOfP4ozBXEydB
hulJJ+qVk2muDHyXvsY+xVE+c3rE0oX5Nr9tHYLspSI35MwEV4zPCftiJPWGdmDNG09TybgQWkhS
CaN7m7Q0ogdSa6KwrswWMtrtS7kU/4w2lsz/vUAU13LJlOmNCuifSmvxNEv/l0nI7B8NHpzL+Kq9
n7SKrUIgNrqMGp+c0VRExtLm22kEYsubhhQLsxpm/GOBld/LfCskb3oEV2ZxrAH7vNVc9jUPM5iS
Q6cGHn80fVds1odcCefE6eXUNmZlzs9rkf5CoSPHZ5HRhuGokUnpiai9XW8YxYE3BM495/HoWbZP
tqBnS2+8XETgtA/uGQjAgDlLLNCGJPIMyiE9+bPshKpNjx3cW0mC8e5gz1CjcpjZfLN2bL8WgDfh
+ZmgE3sepxLpTXVbayZmQY7iAdDQkFCtC6ExccBnevCjhrOWKkfrDzD518DK08QiWXnHqHGFU42d
tvBD2KaIO70BgkoXs2h6kx0wiO1WaSr8s85VneJVL9NqoCwpSpWR/rT7Gn76ZpNCHWcqhbfY6nZ7
6C2CUqXrmkwicVHxkWGa5EGKBhxrEKYa2EZpBnDhpFUFIBgo6KcsYFNAauKFIGdEyYTKW84I/Fh8
l8YRe4tN12Ua3PiPjrLiNSP63CP01ec4f+8V5d20kIV1MvoxQ/pm4Cwvgs9EgeRH0CA570bWsaB+
qa7kTLjo6N82yjdnlq2v/rFCfn2cfQtn3UPPpG1LeThAotxYQtLss13d5vB8CLxKTLdV8et/9TL9
otC+ZZb9BMzNLVwd0cFW1gT/ieUzTzJMUe0NLVxNlzV7O/t6D77xT2hUQ52+BwQVTLYASsD1u5vp
wMLXyy4ZpL/AQQFIGVAYIUTh/n7nUZXNZzN4Vh6FcTwYB2vbIVdTfW8hAhLcS1FT3lIW+Ei1I7Xa
QZLUbSjvfj1BiZ9yGpZdZhSvD6NMe2Su4hAg50qXKjeukA05koPNj09ZS1pImTxbHOpHDmfQF1GN
Oid2SbG7P2dohIDF3YWWInIIxsIcvHkxdL4V1rigDYhUf9pfsURAwlxtHDxUeCTvkYocJbRTWuK7
qobFEThjmsayzD8cUEeTbbgE8DYgeaHd4Y0TxaBCEpvTPk9u87XRLCJWhTZnxGqCwOxUj8ZPxjwX
l7IkIyNIbv4ogBKbmH5N0I3mA4VuZzINw6ZbIPHO0oj6bHHiGo4+E201z/eBDv5Gwx1KbbVb0F65
kEPzYuCnIMmxrrOpJMC/QJvEIv3i4c7ZJPQeVA+qvdbnptb38E7l2IAbxpLsRcroe+QZ4B60ElxH
updk82fR6dPqeLvMWPyz1f8/gZnaX2Ck+bsVfcti9M/P/t4EmSzv2rDE6J1xef7aMsraEb+2Hz1O
h52y9zuIZJj89f0gsTXb7R8+RjOdpVxUY3/FC/42hAErazi3YN1zNzMlOpJ4gYpIySlSKFnhW5Ut
+/hcN9gYANUl1LgVi2HOY+4VD1IwZ8hPzH7YHGhkdm8gMd6Eh+sGU7xhBTbtjibQ1Xt9adII2VTY
C405DFJcZfwRBfbbfGT0ndZfCxkqtQRZ/8VlH5WV+q1NfHtHLY6gsCLEeP81gi6h1As4M0ZaPkkA
7rJDmXn1Fu+AoSPph0AnqGx3wJeeP5G5F4WFHrw8NDsnBdT9RpKfIhi6CBm6IKmJ6Vl50QwZJ9SL
UCrgxLdzhefY/o7xyVQn2dJ0F85+I/YNQXOikxCOKNtKTnsydAn0uw/+F6PEkBuywXUvRQzJwmuX
PgYz1321IthJYQapIN2ht/YelSlahBZN5L48Ob8iHT4fO2ihWhmz4EjiQVT7NDppQRaRhykPxbJ7
ow8CitJow3BdueUm3iGq2eYP+5j0bg5jYNJHb8CmbtRmg/ZYQ5v0ptKOdqcGpjfmcc7SMZyYwUhU
P5eYQncjDbtJxttcRunDHCMZzc7BmHKswxCMjxBJ43w1NbUPwuRITHszenag/7MhVZw4dKSznd+x
ofnaB3k5/kq0HEv2CCbdh6ayHGiwqoiRrUd5zI/8XoVg12c4THtlvvkXWJUTXTy8StsLA5RUu3l/
li7sLY+ebizxOZxF8kcQrPm4ykkvjPaL6ago6+CnJHSLo/qTwq/pD0VVxjQCVNgDQDrd+84Iskd3
H9qxaUMeoX261TIekAOvEgMKalDnwxtqCMCYNXzd2SVMZoFQkwz7erPUYyVmKWCShG4/4XWM5L/4
ApUTlq8Alj343d7xFK1j4fCf6LqvaEmwTt3Y7KfTIqxr552ipGPnnxZW7TB9h/voPJuFF2rZeMqt
6sLfmXfBpGK7/CTCJijqJdtHkNZQkd6+SUmltCTQCRxeNmpky9wwocWDMIi+1jL23ApE9nhCTFc+
rFmMC6Uw6uisBNdsT0Az8XZXvzOHfbZdZmCkSqEGgTslK6j4ufKeIkHBvb/UWG7KPvdJObc9rSoj
Kz1g6rr7ekBjRe0x7qKGL6kqSFBZ9SUKoiVRige/tw8FsV95W/hyis0fIV00dFfYL/5vGHTin3Ss
nUGzYJuwWCg1ldTCHffaylaveeFd8WPtsf/xsIkjp5CJoXq4lGrK6v1t5n5KyDQd8eqvwr5oMpre
jpeO/ZOCTdO943SKpNQBE+x3PljxsvlxXHbrTKD0gj2AxXVWmIGh7o4wk6pDFLJ5Gvol74d+90Wh
4WFyYlxI8nPOMKVluf94buHTMqqZz4nzGYebFMLbtsmUD85hSc9lfrBdt7jxd0iJbD/oBK6UdAiQ
RI/hjso8digk6dNAyATyBAua008eWL1Sx2P4noyGnDgu+qDH+f9UTTmREcMWSLN8JKm9WIOi8uc6
HuXpsslC8cGm4V4DGAqnUz5UDEikjbUe9U7/gp3jjdf4fXKZlgKnAcBSoDStWUZ7xK4YrlZFujAL
AOdBFTbvCsqHAmdSy0IB6SD41KbP8/mu+0XjI2OUhWvhAWRwLJZJ8idSHTuROPq95WjA3+Hsok+C
hf7s2jofsvxuWIx+bL2USHuG4aODYWodNO/ZqQIJU7ijbNCA6Iv3vRTxLmgP9yL2J5J0T71MIkZ9
PfPVpHIvW4TzQXKPuCwIr+4BzuFF+pyIksANP7qdsKXtCBT6iDTZ5twz6bjknc5j17MpkSxed9tN
sqKU60UdYZmf/ccvNyuVIJ0ViK3udLXpcJZTX/RonQqNin5hH1/XMa53xnl17gKsCxqanvcx0XTw
vpOPTxE9aeGe8Sd3Nc3MW5TGSQZBErzdDju7f0Oio1KNb/1EVrSOe5/L5WYd/onXyzyiUMcG+aOq
Dvrp1MvV9xOMDtZpOXdR+ZRYWLj33R8NTH5gh87UUzxRkxR9Z6tCGfamQzeKv+gA2CpfMYMCzV1G
GYmVPxo8recSkVtEW4lZsmHi6POaJph6Dd10zl5q9ZoN+lQh4Pqc5eobrYjJyfkXR5hzjmjnIehH
/KguIKSmsOwy76rYJ74IMWXtWMhl2Y6p9NAN651MiaNC75HrhOQd9PTtM+qGt9+WDADWU6tD1DZD
vR+UdeO8CJtA3soyqPz6awBn/GN9cxFMIUmZhlEPA8AzmPRbDFsXVzqv/1ArBqu3HjBpqCDROHEJ
QW14v8+xxpzGpVR2Odsc0ah/Jm9UX7U2X04HIqT0lRXUyBW4FYQrE2DbzdNRgN1UqSBWL0CrLbAi
az1ehulP+QdwBIHG4aFeEuOmf+oSbPj+8I7vbb6f3PZfbp94pctoKvmbzuWSogFByV2lVjxcO3GG
iA+JvuLZaDrGvf7nAXLu2hpXR0BusT4+qkWue6RZAz54v51sa1WGxR5dqiDBH7P5FFqBNxILKnB1
2JR7s5UMD/eEUzBaonD/wb+gACmPnxFMetP4HREmVAdvVyD1rzK5zgXWzPP/6+kScGGVQKFjJ+Ek
7FPxF61/CLJ1ZgxL7QSQA25TpOaNxMhH81MdnRGrgWUvL6iLw8+eq6s/8sTnFSfQu+dC2IQc1sqf
qIlzmBEkPMmuMy1IzDk2qYQnigkiN9+btByIuBu1MkqJhHOIh6P2cu66E+0lJp6RQ6+Gf/bpuGBR
fXNLqhjtjiXVLqyuDXqwNeH6BkvfkSEnc3V+/wy3bqF1klDXnCZ1qJUMGOJ9Um08Ec9g1sEGVpTv
Hc2zBLPzauDj65KpzjrnTz2s7ABwxHUhlE59yVyfl769IE0zM7tVH8fjwdwRNNr0e0RuCxpWTKNV
zoIDITS/fHY8BfhsbkQdvMz72JIfapjI9VClrRplut1lSeBs4nFkW8kRHnNzLJOIWXUmVe0A2QsO
DgclNgg6MqKtqFzLEikepNhPNjqfCrosLSF2js9Y115rqeXchwkRYyqzDwzxDLHek0gKw0sGN+o4
SKztnKgqUXaOhsoctvIIP5jACj9EVGEiBnKQh6la3gWe+s1X3w03yhHAsULplPeJIHJcptvk+HYe
WhO78pEMqG3eYPA3URseBmg+h/bi3HeubHeOl7U3NmdIaniG9ykyxLs6nQgSc47lPtmg0kfqtlbO
Lm5v5ZgiPQ9fDqDC867pT537Ji3S89J0/3UnM3PbiKwIRIFiGuOBU5mG+LPSfng1UE2ma1IYtsYk
Pr7zmFUANCMJ8I+VCTsorhpodK7/+oy+lqmuE4gmLtCxrikmGRjaXcR9doPUGI5C/BFWt2RnpiqU
AlPTgl6aeJbqsi26KBZi72o8KiEVfOShcHLAbCNnMsbpwVVHz7QPB3LgggmwU0K2k96i7AwT3d27
nQl83VfSQh6TWyqfLUTUwydpyhUr92LrbqtE2NJ2lZ/6HzCYe5gys4yMXMPCNwDw8LMLk6Ym3oYn
hwXBEEFzTvdIvkyi3QabcJMN1FPLg0A9Xmdy0quS76h11ITs3r+Sart/G8hICfv/90ET9UD/VqBM
X0wdlgBRCLnj2znaQKvE1OnMWvoNbRjafyZNVD+9UDFPM3sgaRFRwrvCUlfVHdc+qAGSi0v37mf1
ycu2azY9KZNNXAyxySlkEGzenMqbtYRiU1u9IPO01jbnA0pHU/7PSh5ceaxm9BtGZfDf1jU3Kb9c
0stnZ0vU5LhsmrwpNH+GDEN5tAlw2K4yB8BnVS1g+hILl/nVoD1qLSNxGWykDQGUXildnkdnrZ3q
riuGpVPoza0gdUgkj/9znqGE84f5jrP6lWrSg0rNJuSVnPQ01V7LngPG3pTfv8Ngtk8m+1ZMQTBV
V6Ej0bZ1OeTmQCpR9zJrC3Ba05syv7cuMzz9tGr5ZxyYElpE7algNY5324gsmaDZ0qI3upfUAExJ
SPmO+d2Fu5dsjRh9MQDXCDkJiCs1/s5ys5XlyQ5+6pcS6nxlcetO2CxPPpIfLXTip1oKw12hBrLt
1glCPEmcqp2sxJURFPFyPzE1FkHjXhSJlJ75YukDJs7+ILL8DJbazpGFSLfpsIqOlh10XdG+s3xw
qTuMHV6u9V/Fck5yPM6tpWcy9AJfTnQPv7aWChN+FknNXTh62bVFjykWF/nejQOhh2GJ8iPrIXym
7Ox30ygcj+ChOLbLd/p5Yz+QtwJqjc4TAIOHHfFmYN22JQuQ8oVO9hfKWY6T0Li+TgJBEBNTIRny
URZZWUH72yCDHDBGgYALLAqPnkS2CYyEHhtxpJII5/Uvtk+k4HLssfW5zG3TFrosI0Zcbf9Tg9tc
vn2yu29p+agdc+f/JxiKO0dmsCw8bRiUQN4exaBtcHnHqo9Tj1U+/r2JgLAFUaA7CoiAMuV+JCZZ
ngMiIkP+2DadkrvczXpAuQzo6bifk7YLDDSETs1QZGs3AgvWBhO+FCfCRjsatawhwdz1m6t7/iFD
eT1BZX7aWB+FnHOQ3Ckp1KJSJkNGdNbHx1vfQ5Q2N6S88x4U9ek8I0XZSlhzsJZpb5Jf9KdiIDMH
D5CN5BhOBRy+ktpF22mVDfKQXZXzudd3QqS2c4DLRuAj5m1UMR+TRivQkta9/mllbCAgaesz2JeQ
Yfvm3ztBwPayscHeeH/mIZtrz5T6McVdsMcPIG42nQi5sKotshOXiNMqElMUgdttdCbTlbTqZ5uC
TKoUiuSOpGOFtWt4ST8ZiXZkmbLCCIBYo3XLFXx1td/PimtM1mfYADc6zWpJHgZgpTkd6F7XWXkW
0jFh4BPAKz0Zhz4mLm+L9yO4wTgbzyreY0LdmtAxJls6Jecdgh/K7UazEujiu6rUFihMQ/9NNK8d
fb4syM3GjhBmeOui3Tdpmfs0tWC0pxQdElJzrvhaugqbZvaXGmlJZABUr6VDuPRxFyGWNfsFInEy
yhcXSOu+2jj0h0llGPnmYV9AF5aABNvbAgyXLadSBdXUUb1nthpQXNj3EYCpHuKVDAGxp5JEbNwf
vnOE3Va8GPE+e2eNsd9SmVr6CECMRCQYos8+XNCu4WvCQrv2IPSb1gcCwkydoUBO8C9i+++V7Pzg
CPVmfYvQ/W5bCWY4TscMkzH39EjXF9HUjEftrK9Rfr2r5e/HY7wz/Kh9gUSKcyPM97CqZuITLOzp
WJOYQ0oxph7tuVjy/OjhFPG9N0gp/9HxLyMYb04iq07dk9c/l6VJ881yErH8p6H6/6KdX03IwwTp
4TaH90d+gnaj8WbDPANzKjGLWpMQXHMt59OHtqA3FtqdOVDYGMwXnWKxYuhHhfZ9fJGfi2YoMmXN
B9PaVJcZ3wFXgbTeaf8sUVtmx7fDnARzzx1iY98m5eEdhg74zINeVmCv6dTi6ykOAacLZCHL+gxb
qSRrILv/MfcQ0tDnAFmB4JJ/zh3N0zCUuSzLRYZY7cc3gfHeegJ4Z4FXOGzqAJcHjyrkLaBuUx6o
gN8rXTAVHJNOQAcOyonr15E9zmvaeIzRwB2U9woNq8eL05Ggf2TSXP66huiAqOvEH6Sd9hejCsQW
XeDH18ZeG5UHvI8RVUn0egbauwJ0i3Dq3a2vkl4WhSC/OjZ1aTJmMPwlycqM11ujjwJZKr2eQu6E
kKHilF4DiFaFvhPtmeeOvGppx6OCbcXKxqe59LJdBHYpia1/Rg5hMVQMegEHU3bXRt5vZpn6wjfl
/WDqA4CBZiG9GqQ3aKFPUwrK77OEkhkcQGgF42sOL2UPaRcbMdYE4rFh06VA9xnzrlyva2s9xbi+
Rv6esEH4wR/18Qpe1cWJ6GON6s3QLeOyEQiN5Dt1UKME3K780OzRiMZmPQWitNUlSnArpObgI579
Ox3HTO1Iu+EwZaUuvEwVLWeyNtJShllhiI2ibEk1Wr9d3fbMjsdrlfhVVrAr8S7It5XdfM6CQYRu
XZKaxKWuXfNcw24ZAX6CWMtU4p3N9TIk+iQrGAkw+hUwOLk+dCCFT7lsdLQS0PTScuQN7hi5M05F
EZNha/TfJjga7QcL7flIfjT5lEPE2Hj27wJiydmjYc52wrxD1QhD7UzEOtUkK3N33Qs6jXJhcQoq
SP7BSgL5MzV0MuAyjtrBVo5FyWB3/7Y7x67I9QVYXOFceMAhQF2ju5AmGC0j2QeaAUsrsl1+KdH9
EAgYhHLKJ3CY2dndbqDwBsjtK7Rp3HGp3iCnPuaDnEulRIdAgMaY+W98uLFOwrcdpnwKobNzVUSI
R15OqPTWrfIDmIzprARhXnHvE7kXUlulmCPsDu85OfcQV5GZm1d7sWaKmto9h3Rj7rOWRvtlgqqM
0bbIcX9d2rXIOh9s78qAkczvMayAdwgA1+bqSmOJIKTRity0pFIcaY0QMy8Zk+64Jqsil/rGLfnX
oYMv2MsOa3k/CRswt/qrYPRaBq5+3MnMzt3Eay6UblU6OMhhwq1hngdxQ9Hzn18k81zpKP6oYa8D
bzx/EulON3GHYlKVusNQFI8+BAE6RddRMMJZ11NbhSJoLErCLuqiNUXNaEjjnEZ9DPf5WkDsh0HE
AZhLbo9Cy6Z9SW1b8Tqlva7TBMf0SiUQ084LmBhoKU3iuyWg6yfmA2Kjvf7kTrlGjqtoc6VTcE6S
XoFjEAWrd4PZgQEMbQGzRdEXQrPwrIr3EDLHM8ylB/6EEgBUTtEWyR+BCmv4TZ7yzgluhzDlxHQM
remPyAB5h5jaWr1H1Pmi3uq3s8olBKHFpspvBk+el4HTb0o1Caqtf6447GxvwExalHPE/wux095P
Cpya3TFstCzpRS+OMFKVq5MjZWPGpRGtEXeF57FcyeTqOi1MsYj8GN41rJlupZb46L7YnTggP6+g
l129OsDkaypFTFszz9PLGntUdMxEnkQ6VtLAASY6vClSTgr6CvmT3j3H5ii38DT8JZPsuKkna9Zd
/9fbqBpiT2EE3aX9ml7IU/ULWx+Uy+UUptsil9dBZrV4Ye26OIjQPe5ag8tSTvbcWnKc+tRf+8Nw
Ehb385RdT7rxUD7Lr/e5nmRcQlMY76PDUB5miZk0Kx7J0MPdsJmLTKAYZRVDDTgidm2nQWLqcIFw
jV1Tj8/RiGmIj+C6elqScZACan+pIuE86C9fHNHGvEaF4CG5ea+ochKSO42kZnsP5ezPuPlfZmcV
IQ34ufAzymMK15iSgWryibzcKWb6WjdvsRJlFJNnQJPRLJKBnF/BO/aSsYK4BOKX6YwfUXoJh+/R
f0tUXyg2urH2bSrROPqLbfVbYgYMtBey5FMZ9/n6KDOd+vGBDUWP76vW289FcH0ZEo5CyPzP05KT
ou/D3IJzUFaH7JwHJqzYN4Qs42+zpdfIfpyWtnnwgZetbBXm0mJBZH9yehuXV20DxO01KdzYI5/c
glo0XBNaCC7QHv8mKq4HBPylSzO+gVBtCpLw/4fv+qixUwu4De2x2l0ak49Ip0v7FGYWrpde9pQ8
58HnddvEMzLTTHF4E5I+xJnNVad8nrECY00pen98JlMHb2c1YHLu8Le9LdTA4NoCTp+9iK2mswg5
/7H81SdWcrWyd9emEMIwxrvYWTs1nIezrrFtqdrvSutElriZWHUxtBG4I42s9t4GYzHZ5ZYb/+t5
WZUctbDhEBjZqhbIgyCa+pLt8S7bCTzBqht9Mr4MYtOEOK2v4pwN0dhU45VwCw/3NRDpEjt56rzP
buMUA4LvbW0L4UxCSdLc/Z/kOay6SUU1LDGLXWvz2meUulLD1s7RLdgyPe8HFHzrqSyhFCjMGm65
5pWiZpQjriGTEO47oLkDHOoIUS+Y4lergbJP1A7h4/rryTnmudDxJP1tG4mqgI3hkGqHW7uMz6oA
F2YPFwtS7+jBoOo7Fzn0u0BPwc+vbKNBLkRD3IPzHCJ2DBb15W2v5uz8gqO2MKYQU200bfVwH2eD
VL9fAQ3FvMq6hg4MQRQ0WvF3qs7QI1LMPJAM3FS8M1ELFfvEES+DAS/xCEYuRkMlS1RQmbNEu2+2
g29CjTSvm5vJp9+alAR64YB68RxQQLiLeAxfjISnYyagmZHT+lVgJ9IT4NXyb6RM7yepdYGFpLJj
BnKhHoB1hMY64VkNMMAkGik9SDqYrvuTBYWt/1+oRgbyKAUYnbqWbwxp58KvNXptvdhkAEKHQf+f
LdYKSrl2NSgj2HNO3Fd+/H20ewNsGNJGPgfySfRdrktcrBVkSCCJuShPxFYJpb5Qo458KS1E9l4F
i439aVmfcHVWC/liu8OV7ufdF42e0bSngsl/DryWdKy12p6BJwWh5vgdnvK1ElRqjpS2Gl4JfqP+
pKwJ5U1Brpkstg1+mYJMKnA0T1Q2o5a1mLUP2aXWn64ydpnWfsxnLoAUc1tZR6QhbFAZdoPFPCk1
LNPRLaG5dxrUG4sbTMR8G9kM/H6exFYgWqLuq7+hdyuv2wXKw+NvgKM1D75o6aCrpaNk5iWM+h5f
/vJt6ko5AeXzgrDCK4KWSU6BzeSP/+J4uZ9KVk2GdrLCrWAzM818TSPmfg2K1zFp6ljeylfnBYip
Y3nmRKoYTaPL8gvdy6djAYa0DrDR8j5a9FqO7IQvJoGFekC+tmuVUF1MWOUfIufQXDLCHyxlTtBA
B/P5rDBZF7XwnYgN2hSokhhAXf7bTROlUHkuowhW42LGib2CZitcRfJYeef6Pbfu2DV9idf5p5n1
EHquU9okWb0HQ4bOcG04rbpsmFXjzzHuWSuEXfj7t1T3Cbphc9g+9CXHNJeW6HMLspdPwGc3Lfpf
ToJXO9Bmvf3yrwRGsvpmk52sP1oLiLZcP1brxih86WTl3S+g6lrVlJl5z4FBIaUFtKPCdXSQivGO
3GSXD10pf9i9EzqB19YvPFlB5v75sXjbe5CehPkioZE0jVX0fOqqfZdHnsJ6aq/0IFrFq4l72r9Y
SqiIa58/ljVrb8mld0JGAgxQ3/d/Tuw2rAylLJFd9EyDCVWph32aw7nmxSWcO+RfB0VCnalpCnIG
ljFQrLQjHxznsrIEQWTYf+t2AsEwDjGUsVOGfnBXAfscKxtAPYjjgklP5bXSarKnynNS5X8VoYO9
7xurKI5NMPG84DuoGHzJfff+HAKNzUEagk2wkUl5KjfsDHNyddNulOValkZfQktpjxVP3J9jp1Uw
QyX0p7A5J8fmhTzHkPzf4kV/bYVBBOfJuBdBzXzab7FyfDEymUIRq02H5tXKzt4GDFfJxvGqaeDJ
JnNlfLsn/Vtb9qFwKmUxorELYnjM4hOlNC68P48SnjdmV7+T+s5McXKfkubz4xkjaWQyWTjSOhv5
F2RTkTNDSurXOn4lL6HBoPodBTKqqsqM9ah1LNLGENevb0f5Wz5x/n5UPjtyaRnOGTXDaOtjQJB7
1K5FzA/UYTcaE59TCk+cOu4QpwNgyu83UpaW8ENRkKRdyYq+Va+PYbl/pwH3zZ8sbP40LiNUr8/x
u71p0r7hZlQLipxcfkgMZEC72he687ucGB0j8/EKlueqQoTS87esnbR+2FWpAaYkwzMu7aVZJe8W
0fHsuipeJgQ+13sPnLqYj+YmdAIzQB3DlXTCXUKG5s7B33sHHF+SgP3M2OhrSE6dUbAzce/S2CjO
dHhGAqmj6CNHGRTvnYXbnd4q5OvOOQFmNooUVZwZAKefkyjqxlGLBo+Kyw2dZoMlRLOjGCQX71IN
ZhcaJyFNdelNytQfs3zmRfEWPnHKlSUYOGkyOswHtxm0toP4i95g4huGGNhjiiEIT3g1bUunwUQ9
MR8IjNPZJ+KOh02WDPqog8hXDORQrcZHeWmQwLKpSdq7NbpAYp4ZsTCXR4fb2sxi5uPFiCjiCT1w
gZNNEXpxVFJiBSIScz7RoEMCpJUm7JU4kQ2DHx5cN/IsIXgkpJ6mCgcjTVuFQpVSgE/qcQbhiy+0
OO+1LYvSXqCnSAdJJAkqWwLBxpBwtRPRMKH5J3A8ENIOG12z9mA5q05GQJjmHx8GU6GiLIZJHH+K
6ppob76od8Bke1CQf1TCjg/FdaWuJuSzd69au/ySyyTdjMOhIL9USxdIbj5iBUTsD02Z9Bxlwiox
MHDSzN4Yon7olaAkNXi6+s6Anu6t+ZU648x28bb8hzIh3Ny/gPYdKhZKie8gPwR2jHXKFI1icS4I
DMW19kGY1kdoleX4JZDqVwfRPVGPFUJrLpP1xtOl6g4fE89FK3yfOtjsF/q0/SgogMG0DxaAB2GV
2HtLdt79/dLA5nDvIc4xTl3n8/q+DLv4tYM2K0goGuNiQS//5eCS9rPydNkt6jQNuJL1AKLx2uKM
/HWJRGovijmGjUZV5+arrcqt9g3W4eKy5av1eADac52PGB/n/x1g4cH4VaboFjPQJ0Bj67NWeS5X
hWOSKfF+igbo7415j12d/82cY/3dCfkpftpV/5QWpfR9dPrrjMqzkydEaVV1h48kt+PhfFXtugXY
TippPfA5sUjQa4xXwCNEw8anjl7uBL8bf5aTg+C8l1ZtrJdmuHYTXCEv71TEDC4Np4smCExB96Gn
neNvcRJfKst45ypGMdeUrOq2ZSattuLsLVzD1xhdNmsVujsv+ZNRxCJKNkH7JM0uscR433C9zLSZ
a3mtUXtxkIO57D9kJpHkQL8WprhehC7skvXVEuXcTAlm8Mw/nXf+BTzeAyOq323B+Zkhys3jOplI
Z34J6xdKojfZWHoChWCKGkayf+SMxbq/+5xKn2AYybVHpCTIf7L6h14H+TJq752DmNiH5NuyISeO
JtRXSk4zkuYpgOiGhyFR3YDIPH9sIEi4l+vJzig/jG6qgoD/cEEpwY6m8W/QeNFICeLgF/9oES0K
TH1SlkM57jZdGMkB0oKbhSNVQvknVhi8EwRVj08rvJeiXCCYAiGto2p6ocPhbW6iSNAS001RpXOh
i4rbe+XysC2ipzIDlCMARrBGdT86S0KhmeMRO2ZvM3PxOosGzrAhViAVQA0GMjClRU/+eHgeaamw
KGFa5XbCKLqatLcqZV1Xv1wwLDSxC6uQ3M87yShhzigC2dfcl3533c0Wt3HeAKXutZBKHUbwBKaG
l2oDlD8xdHSXwEGsB/3YkkMTPjBby8hEZ4HsPlmsjZqERVeZZj0wuU8WDvqfsNzxGOiuYeVfYOEk
ro4gFsA2fV/NXRx50MzXMZ6cGWcJnKQaj9woMeranN64LqzfAXw5l02xJXMXFXh47dzU8jHMjIVL
WEclMkWMkBZNE9Gi7cG2cESSf0W4luxPiwAQ34b9/EhYXIm5EiRrbUBgvaWlMdyVzjvghi926duI
IQfY/JqsAy81KQmmRJIETcsII5yQGIIlyNj07u5SWf26C03GPpgEf/DW0CF9AqVmv3XpQtAivyjD
EC0/h21ONm4iAlNfETMRoBOlltRnJ1xD32JWHeHA2APd8r2chriUqLE3wEVMiDjnP3t2zGpANVdp
FGt+zcZ0va8OvrUJWz8q7SU10LMRYxVbRCGCyfrYS5RS/SCxQY9XUACz6YxXv7338qc6bNQwRTwO
ClNkk1Np3YBAl3onlY22oEA4Yxb7D+3VlN+qIQd3lNPeyqjDHFQRn3NIVtKjLBZJGLCWZkMcswlz
xI5JFrqF5SKI8g7bFtvdlF88RDAM2IViF2jN/It7KDu0ISW/bsGtDYWaivkS4AHUV7zDJxt/SCCV
X8m5Yx3UaUCtBnfdUjO8XFRokMpW9hK8cmFxuFlc1Wxf4LXiMDZowmIHoeF2QNGViIAlH0hxj7ca
3T1N8rFYV5fO5ZRNxh/s2ntpCyO7WljAs11QqsZ8ToxQSzVGm2xzmjG4lxOQFALcZltjVOdvjcO1
ReSHIoM17aOm9CBcAcuNhvWld/QpUdmJAbuqoLYLxoTf3P4LaaxDMwkJPKYKcDj2dzenPhKP0MLq
jh27zOscZAuO3Y6Mr1DqyVpi45Nhnz8xiM5YXZj3fGeXW+PKJR7t6kjiTY2k0Kwks1LFFzcbG8br
dB4oUdf3tF0Y8Ds06WfiqeGyFfPhoe+8tVaNmq4iUcVK2ZOw0CIZstrwRPvnbCccWbsiOw2KJoMd
28DLoEAuFGCIl2/swuwUoXZZwGn7XPwpoxigaW2ZkaBOFdr80TD36g2WVHkDhzGnD0wyhL4P6t8t
jH+56lXbUfKDhX21fgKdOjEkO2n29ObVtTsZGQnl41BzsB4mrmMScOKFDnRQWKMu4ncB9zX2GKFR
xSjjB7vSAxHplBv0hImGH/fu66QRVtrvZo/CQdYkl/juJa3XX04omWE/trMB46AyPDvpa/Xrhl4O
d6ugJEwACHGeg0VrKIaMVENYX9SB/k8fNVVR9Js3fTvW6Gh9cxUebgG6zkxAyYOvWr7346RmubHA
H3RXUyxDnQgMgyZboN908UHys8DMEGN3XYR41WlnwXT6pO4pNF40m+klIhBJub2Sdftx5aJAsLG3
9Syboz2mNowYPJP3UOQ6pisMA1nFXUId5o7XjUW8ukfy07aIB/Ar2fAG6gJKFKDgLE+O2YI6nhKj
UKKVT095ENYG89fisrw9nEzBQYl9zsGboUAihJTWIad80l8XMcIXE+Vnug4XwYZ1aDw9XuzCHfh8
a3yWm6W7YmHfBeaCTSB8z1DOWmSDDCmhx4AVTyB57siR017XFrMS65DaA7S8w7hzSiF92hZIcQA9
hkhQ3w3BA55Op+pjH1JXm7eGgrWZf6snsLjPZNDSsV9IxycMrRD1Qy0l8F7coVCyFNKYaVrWqA4s
8GTG7jJfCyVvL4JQ7e4iKDS2CPxPNlc+M69+VDHWNoVWGU36R9z3KldWar/fftJlTthJrdd9Md4b
fjHog5qAXZgozB2J12FpO+FaI1+2jxVyMah2atf8mDGSQtTKU0ZrLzYVPCwwv0oH/j7rrKjVAL3N
chg9I3Rgrer8kKqRRdXZF72YQUsdVsoKtlf/He2gZqhmZ0z+NX5lMUkZ4MyIx6L61LjXVw3RhNax
Sir7zi3fM/yrlBOP4tx66EKx3Ez9oqSb/VkAYnRVsbLxFIbeiC7GRFMKzAbalE6nwULqkQvFPm1U
8r+lf0E2ufrvRRnQwuQEtaBgp3OwgLMFw5P7oHAajtMpRbeGwtSf9ZyBvmwHq1ubuUoqIIhDDEcT
8QX2dKoCWO+JGgNfH1TRuVXXEUo6ZawFVPlitPUP4ZeAtGNDlbN0D81p/cMsVxwym4KBNERgNrEJ
DqbBcOU11mOJLTiti2vBHWBm/EtWgVwhrahr3V/ubuA2fixYBxZqwn83iSwZqfFUH+jdvypItz+0
woX3qzpgOZApxCO7UhZD3/teDWxSJ1NaDX3msrN8z7Kw/66b3FqBo1hgUS/w3nXdLd1/yACm1m9y
rbnQpjdbGHNnHGVvdwGqtxoIrqm0xR4XYPcCVqFHHSNBv5b6ohBJY2yRu8p+l/38D0U2tWVFPj/v
7hBOZteNvxK6iUccW0IPtMPvwmqYHkLqYPPE/sahwZIAhF3iQnD4eFv/v2sv61ckwalSu7VJZKOH
6GR51uuDsy5HoBxLhm4PWpwb07ow6IfLyyPVN/h92FDjzh2CWvBrQQ2eq2Id/72/wXmlclegwB9L
cAGoFEtPDlvtofDtitJuN3SsDd6kJMM0iJIrdsVokBEyWUQJtTwxc6qjglwV+nIhONIORTGMqDUN
fpg7jIc3xsJV6osQXLHzSD9nN1rUcw/kspuOqv4XDdxMZk4e4XTLFb1mmFDAJsNHS9k0N1KswoYY
WCx1lPhEPu5sHjH4u5SYcXzG9kgPbiFBHt9QEfYTI43RsU8d3AAr1C9JzPuqLjwKgYVHr5T0FnG5
9AP3wjqjovl1gOouWBATKQGhiZpwXvHB2ETAA52NBRZIDiqhttyqtGzKgekvuoo/RORoopeJCeNk
OhlQ0dtrpkcJq3/nStVRN/Cs1fEtl5IlOBFbc5ao/ALnOnMXgzXYkPCMNI2EnJ9tMkSsfjVFqQ1I
oAozCiPmH++uJmXAoHylBXSWfOZnqkJPnfY6jx3O7laqk0/Vor3p0PfjMp9h7q+uUxzms+qbozTs
g30P6XFCyQ9bA4CCuihxzl8AK4h/RUvlFMXb6PQE+xPePaxdFtousEds3vDkIGqk9MpPlLgNYDF3
AoqPydlYYBdJkYCQR3uXkPHL5JYgBTwQu+egO0BBUmebRihizvL1lsnLyCafdQ2YWTeD37vFtAd0
dcSV+AcLuuAg8YqS7964TcPiuWxVcvampcvsfJZV0ZINib/K2eAC++lWBMmGm5nIDoBaBDK4NxcD
jc0uEfKi6fElyr5aNGH5fUGGgYCRenUKKQ72/CVkYUGePZp+lNtJy0PcyGiIspuLrfeBHhYrfy9A
9JlyTafn/HJsKfGkPTSgaCL+2wp4MFtRv2mQcVk53mFjZPquu/PnaFvj1Knw9PBnvMtSD9eT41Gp
U/eHivMQp8SiHE/kHUY6IW21WnTrlFIr45O8wOaWRKEzxfT9IqFic6Qak7Wg7wsem3vDflkbzYRR
1VV7nTjJf5b3y6fEagXam6GtaNNnTaFlaIZ2lKf9dLaou/sOQ/QVVDBAiVY2HgZdan8hoYflELUQ
BdMhUqfgaZFWZ1EM19uQzWi3U0Qwp3jU1eo5Jj02s/0eU30vDL1a0Cgb+ah60Gkztdc7wwrwm3Xl
jG9jjj+QUDzFqFqTrqx6ZMb518yuvZSNT6P7T/E6pg5tInoY0zJwD/P7kkuL/Pfwo5UAGQEQFBu8
gXM7qc5S6J3Fg8JPXSeCJ5m+7jB08Lx2F/CnGicceHD+kOcGQrN93CUR23eKzspbCT4QvHhmUXWo
D++L1TqPzBMsedR+SUqRIHZiaxPXskPmCg1b9wkZ4E2ySs/hWN/3hDvULztpTWQf7sUQs8Z+xQDz
vHwackpaq8H0ICRJFbqO2el7lh+DHwQrqHyNx+DYGW5t8/f1i6vlnzRVaksW5+fWWRPW4uAYso/4
P8JlKrFK/JDUylrG0VbyaEZA3Rk7ClKlV2zlYLHhgz8yDVFG9rooFu2G+EMy/aMbKMeM3+Cr0C4x
279D2idZOVx0rd/0HtmdZ3cGFjHS82/XOVp44KII4NNDCYVgd5Q5LMkTgl1KK6YFgDzEex3coN1Q
jBI/BjjsL5nOXJHpRy677NuHIQfm1Rtt2aYD0kmTHewPWImaVABH/3RJm5EnRlFatQypf+oFLFLE
THIKNK7KLpFZfF5DknBZi0ngAdgUGR3GDSKQsEFp8bi9viSy6xsO4RQxtfLoJBAco4Kxm2U0CZus
xPg9Q/YS873iFOZf2ZZitR3o+OFsG5/7Adejr98QtRnYbK63BtJaaxQlxCLOGkUWq1IvC69t77la
zsTZsnCgqiya/oQQnI+v0uydYGIeRcpWyNDgtjDKhWdUuFd0Cuc9sXRV8cG8/FTz4t7lq/BmiON0
NU0GV/uKUoGOkxm44BKXtzd6RNy8w5pQOEeINv9A+ZsjQbGTdcxAAiDL5wXlS8xyHR0UOt+DEBbg
7Diu/9208pGs7egMRKbQA7lcTEQgJcymSEKY6k8PYSHYgMtE8oxCT0879YdIEFlWTAXhQ20BWH6k
YHAkyxcs6ir2FATqyDnq+Z+HHQ/bt8dhJnXTKUmeix9wz0zEP116lywzasYDmlbyh0oVOdbr/uOq
YfjTvRLSQbObUkp+dk7NMfPi0si/kYtEqXxW7/vMCWf0ByNip0c+oYnHwveBq0MrTb8odoumVv9X
xd299wojXxEIbsyQPKd961TdwozMr2cxYcFrthewSPHFDdh8H0TYTTok+0pKOhRUH+ahfbD73UWD
TKtNlkmDO1c12CIVIsySN/Cy/oUaonnWobnuyiajoCCrUPp2jtH0zke6r4s1LAhRUwRG88DgW7/0
7C1DSfMPnjqfpr5cz2tOwpdxcp9pfi8ghpF3Gf9ZHNIigDndZDbJ4JblnNNosf4NAlU1CuRKSzhu
1FRs17c1SbNC1e5g7mo/1FnDUrCLw3nLOcRL4UyaRCEL1Wd6/mGMLIGMQgjaBYNBWcWgUU/KBaqR
vPKK+Nt7OubVprd8WCdetEZaBM+/3pT+0CYgZslNPRXVW0ZeFHJDPdMQQ0gmalYEDXrnD6LgqLgy
L5JpfOsCZxq5NiA6tKtFe6uYp/MTi2fNvfgcLf35z18yIPiIaQws2bJPvS1IcM5yAQzGE4+oJjK2
pbLpZDVspISsAd2X4UnJJEsMnbsjv8//SlDLbCWYxeAl5VHpwEztx7m5gY63A2E4yMvS0F4N6B5L
ZRG8bzgfXlSSI5Rex8nLcXbvHjQbaUbU5+/oQ8wKhgWZ5LOVVZn03zLBjX9W4jIAldJWeHjIO98q
AFHgQdjxgpN+EF3d7UvwVJ2ktFEGWt1fhZTRMNPkNS/SuhPTuwuwuxiK13l3uUP/VMKD26QP6XFH
xXCDEAao7a55m3Ca8Ddr3ICbTi+EXuIWRQkbw/HbB70+xQhMLvXVscLmt0HBD0+/2wsKAkG0j6MI
9Kp09XVd6LtjhvQe5XfJpbEVzbkFEBTmIyf3kVEifb6kxGMQMcYErUYLax3oyd4H9rcmYGwdPERJ
SupWRXW1nlcgdr6Kkb7qDNJxPfbpDQccBsvr04JtQgQdb+1RAh+VhmT9tFNidLaohIVGE1gHvPnw
IdFXVdgtrdRJmff18RJQfFYHmB0eb4T7oFk6t+lFPvdYBzSrlLWJbYz/pRoUMbZU6UwFHIayrPps
nHt0vgpHkhI5o/czk4WFkZhZH3Vi1xizmGSFVrz+LVZu0yiu3Nqv0r50k35Hj2DBIcacp//zuclv
tXinaIk8izZZuDG8RR+TutLGJLcLNNU+ItQgrUS7MLasETkTkkYKXaBGz7JC6TucApQEkobRn0Ru
fskOFAdPwY0MVic13JLVLJjFs1HqrO5hVQufBdSvqjkRuUuEbC3SCl+1v5ptuwU/Ei3HD66NK7LL
kJ3zuyiCXVFc7D40ZLW3zLOPCIAiGz9BfT9m5+eKozPeuGgLroGsPCAOmHGcE8A2KVcmxb/QmYlY
FGvivG3qVbiPYwplgAny2C6XRxTZRzsjAXtGjLYAoQD4wu4BBNesyMAJXRebLInSsHpygpfFc8i2
uI4z1v5yttgFpXGgM/otJfmf7Grne2DfcRZJ5TgKWAVwSUOmKyAyJh445dWxPzouu52aFsp79LpY
LRZHUeVt0SAzRX9wwgOdsxycuJLYR6yMsJBF1v73mA13CG0wZM5ZBBp2fpbrgY5MCItW4KNkyggc
Q/fTuXSSHmREnFhU5Qbn9hDfNbHj/wgykWYIV8Chbb/ckCH74MkvmWA5OXrQ2DXnNYhvSOcHOQql
zHbafmqGWLladVqiaxy2vJS5HiyNfmzr/f+LzU0PX05iDMt500R52Q06MWiWIUpXXC6CR15BncLh
SBoqiuOVu8fIQtsdYUZe7wRiIG00ZULbDK1W5jHgLuIQ86i+Zsmp6NHOIXSf5cKT01MnkULTkNtJ
88c59i/aVU4N5zIU6g5y6Q6fEn8vNdN5Z5rHWMMCraLNkP3A9RQLUUUWnznKGqoDh0qlWuDN4dPc
rxa/fEfqI6R5wyAz/z+qC45GlOuRdtXwF0K39emQWoFwCKZpxyQQsbCbXctU3k9JAiO9Uq5518fl
K5cYV1/X2z6poX7Pqy8kDJxY/VswEV7ggGynaRu/QSoGUV/OaRUhCnT339VJe3XZM2OYMmJfPp/+
sOxIeeIL9oj9ffOzQ3k1oFTjcjMNji/jySPNjYeEImFGHSbJx7U3Sq3PJ7TPhgaA9a0WZj02EJRG
JK4XjPu0cFdlhPy53XQmgHq6aMRFUyYQlKsEuFbs5muLvbsVh7u7X6sNAWwVYaH/vKtnsMPgfGtX
wKAzw2qdCQupUryxJ49gCWtn8ekfpSf9r8xH48V+9A4GIDsvgZ2UE3qUU9g3Ua5DprRhoUzDlLbn
7urM2s6ea0ofsm2n0zbZRs4a1IJTV/1BPszxMpYYXqXz5XIeDkEudPBBB7+X0A+40ldV10ChGEJw
TmeZfXinh7Q7OtgdshoKxlGsA3jr5cSbvk4xrZ5ljisifw/VgTC5OLv0suKU2eMM1WsWNR3MxYjy
7P6LhLYiZsWChPe0Ut/kABJrHqGS5ZrJVi8094CJyQBYq0WLit8wu3Zqb8giWbjX2dulOFdWS2X3
aykWVVbGphh8gPY7KWYROdsyoZKPfeP3MD0FgITt6LW7BeTM4DkQEqciCnptQ34tVjYvw0nAZ8LW
Cf4xuiKRkSUQxSnVB4lZkBhpfZrX5Q/n03UZLKuz32VHLtxWYHHi4as4XoMR7bwz5k+DDLkPJHwI
gq+tNIihKIjANI6lmwP33iBYRkicmLSR6Dv+lyvXVaFUgkLZLU1lNk5Txiiixe9Fs0SF3JnFkQ7K
m3CpQxfH1K7cAESYQbzJYNcP2myGu/pAig1qRUWkRcm5wyNv072ki9B8IKFVU9NyO4fjGTzlsDDR
9EuKaHT1gW++XRJFvh/Zm3Bfl8/a9OU83QHmhCkux+6xrHCsNdmx7n/w6AS7AgwB8pViRx2HK/sM
p3qv3SAeuAS2mKFT/o0DrRdQfducZFi3seeDoe0nl2Rin/WVdMz3SKcLUJMAr6xzE5KF1xkYp8GV
aiEfgmXeAXJySA0OmbOxt2vrzosqm0ZR62LLdy4+Ec+bK1+wxRTfchYsrCw0rKWFev1JDNZsT1jL
NT81ieSw9ym/pKGY6wDdeND3S9Sp/iNk4sKyY7ZdYjO7wZO1g2fMTpevTPbffSEjawTalHFwfzNV
zGkhyTprTh2w977jekrbPDZ6kM5QEbaE+4syVg8hiJ07Ie0Wcgsjfo8YiO0S9jEorDTaDeZ9mHdG
tKy66Hc0fr7+R83rprPzoiNt/DLeJL9TGeUluT/rXn2vHDeL8DiJKd4wPlrd9TdSXNvw6x9yUBt6
24VTI538CYszt1/sM5ds7UikeDSKzqivrKRuj7lmEikyQHZCrLEIZKdpKdCG003TzFLL7Ee7JkWV
iFtIJl3F2UXEy/dssx6TJBRvILJNXOJQk2coVvaPIrx0m5OurWITw0MSI03r7zpJnjn4iRxZCagm
bMck7gKGIFz7QZmfiAyWl97mK0Nwj6wrpMUg5xRT3tI4uFTPyv/VBXJqfQbog4xBc6FhDGbNWr8O
rGinoHjNv4fPFkPtatpyyp6WUMDp5tUmtoB6RTtahMb24do8vTq9MEASIU2H0O6CMRpBLDtlRB/O
J1SZeFZmyix8Y149IiVACNpgQP/7I0Bqysqq3c1LpbUcFs/5fuCdFc4D8i9APoSrR+5pFt7WFYYL
Eq2M1Ft0TUL69Z1w5bXR0vUqC3ORPqv+5gQNWMPkOcFrA6prBnAAdnsI+C3BFLuQZvVHeObqX4Ow
ekU/U1RWyhpEpVzKQtLeiiX4nqaZ2k1XCGJBOAwHP5F/tll3GUJ/Lbmxw6L5qbA3z88aIwomjm1/
CQ95fMhuLyWtXevxhq6YI2DLhsgnke6jHiV/qWddlvYob/yBUB5DmWjx4Ne2bWVKEyUONg8PgTVD
97gb+GXNoJ7Kq5ybrhYmv09m0yycZt94aGNkGz83Pg2zQ5Mq7RbAOzgdjuO0/3c7ig0DWL5S1Bf8
Pgvu464k2UFM7A6Mp9V0qY3+s4x9Pe8yZKeUp73t3afpgYbR5/w0spiF3n9lwj4SU12C4NWXYliu
9VoTsPLynIT3+id+x+iyq4bGfKaEmyFqswXTA+v4fdfUEsvV26dvGOkM1C50hWno58yecLs44lic
DsenYeHsKLQ3gpeKzVY68SXJj7yhQjSePegtX/N9BksIXfIV5w5d9g/Pvr7AAYunzJ3UvQ/uAocn
K9Jcfxp+hQnzauZEVPXNtrQB0kJoFE2SF0+Fr6uJnqPyTTmr+QQ3XXrjxrzYXEdxREX2Z9mF/mpm
EUYfGdWmkZffCAu4/p1ASwWlsw90yU+xlSjaHgL+m+IbtcEsd5hfFbLpHOUIXhtXeyuHQtS8dyAn
BQ9nWnBmtVlSr/ehFbFot9zUCEz4eBNuJhzSTIFFUgp9mud60RFXvHc3cVpWRLzxEiQlt8dhDJ9v
FpwUN5Tb3ekvouzhGrOEsCxmdZftjRXVMVNehgpm9Pqc+pl0eeI9LdtQ+hRCagot8mIF5nC20pZg
qbWlKjjN6s3iFpt1yONCzjJU53CPLIvnVOarEAjx2boGjWKviJqGl2at/nW3c1mbmJJVeoEQXQdY
kZjRq26/NoQjTrIfgf5OsAx6W8dhyE8tD/JkjZrzW0f8qUjulZ8EC+LFGswtwhAgtTh+I3Ryavzg
z6wqJFjvfRsTpnk+LUq43YV8vN7wGbhUP1ibIlFl48QVfmkhcfmAUaUJUbNeU1EIfjrnRgBPcqAe
GE0QLL6f/MpK4EI4j7582lB5d8MSUTCOO0xT38evuzaTEQjU/h+N23iKGKpACGSyy2wBnsud/oxO
8Q8vIhLX53/4v7uusbWSa7LQO88RoFb9UiHTZi6MZ0xTlGjXJ6AY/L2AyK+6ppP5Wp5BGclNAUar
9tFDBfUFlxWmWnEKeYT174ib+Tb9qYG8YEo7WfVsZ06CLqtVGb5qqsk0Qu9UQfkPMFh4E+i2f7IL
RHFXWm14GfL4vCl7mdKhsuN/bjrfsL0gM33FS55il6s6+wzWNENaUtUL8E2FIXGfRP93ZAV3B3mr
IV79E7jXTtIl3LxXsK7YdRMle+8IRB2serzaUhz5Bna2rSdRfyhUQT6k+3yvtIduOR2xWlV8kqZ5
wIls+BpxrsaisGlIcfcNJBCp2NuuXX3upeIc7mUhKbUCkYAztcwDJsq7tifd4M24nhFCFeNjqB9s
70JyqLrNtEGgzhxZbp7W8szLQsBCNTD3Nimn/MP6/QZ9Y0hhJ3biqk3RZim/g+hv58Sr/6LBy4rV
ZVqEa3bpHfLQDnYeTWWTBmu3I1Pvq87d/roC70PSNA8co7ySmowj+SKZmQ82X4zxnrBYeuBOf6S3
3ARML/WQtg/GiKG/oQe6RO83wcsv1r/0XI5FjvDN0VgDflnhos7y7Ab9ALd3y4DjJpkJFgMRXo85
SdUMlxNRwz1GyFCOe3ij6emAxQq+bW2/SMQHUkd8eeomyhG68DPOC1wMBsrtE1YISJH0fi9exNXT
kfg97peIukfJhH4B6upctr3eq7HLuoOMaXF1tetiFB/9m81Ew1vqlSsyH4MPvuq1nb7fl76PklQS
YVcU0ExLKNbNpx4CtDG00mopib8ZE3SOAdW86aiZUMg4nZ/IT8QrvFdm0E9XG+bn7VNHz7h45ocL
l2LZU4U6xVcav+gs+X0z/0/td6k1etJfqqDhcW+O4qkArQ1OVqYhQmGaFCy2yBNX6JAm/aypEtaA
V2V3uRhbGCGoyc/ZYtISeFtk3Gl1F1b7guaxK6CZibMjt0CFWX23N0yGAOc8C6d4EADCLojfbMVl
vDQ/2q+tA8udVDgzWowM0D7vLs6JLzvJ5CxFA6SZ6G6smtN/n5iQuAWv8kIUmqeKW1fzj+N8f//6
HNg80x47H/v51Ozou5oiDiy0vKN86MtdI8WeISXfWugF1T0EOhELqiivMBTCxFZjxtuAa681MAcM
9pVdhyMhE24jmYcdcF0uHirwxfH/jHFg9Eom0nkT9WBuXYVTVkfQyN40wU7rC7agb9Qrtvp8eJ2J
yghGEM35u/NlHBFNjZHpQEcF/vsP4umG9mUWvKGXybW8yNEBFeVW4R2xvnbS0ZrglESsTLSRE2EW
LCLFBJDAb6J2HU403C//ZgrPD76Wka6HexYwjr9TJoD5Kc0cXJ/rvV/UpNVMeP6TcWBDwW0SMOPT
ZRXHeXd7GQK7i+LbBtfcFZ8NfTaUv0gA4UJIGbepaSwMd/56S1+fwNJPk5iBu3lFiCIS52c3bo10
9S6DqYA7gFOYglrBf/JMyk26+5tY1Z6BhXi0E5cz5D7Wu0dG3zpqXZaJs4Y/hPrttU7pkLznX7DY
PCS/okXoIQhzc0ZB97uT6yHDP6GIaFNNCSVIVlTz+lk1Ru0ouKeMPoGe1Uvc1gRhlZcaYeKJyMOY
6CKzZGArXXoqYe1o9kSMO03I6jTJvl1MxnUPZR53QpL33FiQJfZxNMPsMR1I5lEsJSILGcOZGXUn
1508IAQUoPqfnTDrxWnrMPlATjWUkLpjtqdoPe/1klaPAtiXCPEet4ETQcNXwFs/V33lVAy4J8Jz
3LoFwtXb8tiGohY0EabGsWisb0Vks0psNSxL1VwdEhjLh8RqASUoBFUJ5WrsWu9qulacgQqvvu9R
LT/4GL9P9PFl7UbwPo33+HGSIPAoLNaysfeutn+GD3KMP/jncu/w4+m3gzqMXHvmETjir0M5Bln6
yYuDHuBLDQndXbAQKxv1khGgSpyUTAoyTnd7TfDShemG2HrAMp08sN25CCM59j4NRMtRSqPAFMKQ
DotKNNriQpAdt9GO2wiazpN/ucI/y8JmwYeD6iqLcZHXvQ8cJKoBz9732d8nHNP0FNw7TdUMWPAH
fRIPAfOQ3GuTFCrYPAZXHxQmroCsvY2Mw3dRFkSGx55qODTZ6kW5/9TefPS4JKRdCcHsGWrEXqRA
E2AfUeyJfdaCPK+p7XVIISXL4ZlASsqTDF6haE1WliIUnYiPXwykWcqVoDY7qFJoEYsgkmHRUAcB
q6OSF6CAfBKO5FX5UVgjdPc+oWU4eenoDka4LBTdgYaIb45MSBPRKk4kPj5EZNwwIFPtwLQilUKG
wPzcBEuJ4/h7q+XEsRZNxSQrgESC57ltHFddKbjXrIhnUU/A6VHdqUo+zDCaLaqsm5uQyNzNmAMx
DWJqpfOUqaXOJ3b+b8wtoNHVrnnCJKWUjQrQS6rVWxTr5Ps3LLqE/tFvU1lmfsF8vNcCDOMzaUon
Nu0SZAJAj8eUPYFVJBCc2S13smvRmfdozdwsZR64O2xHZIf5j7X6qe28HHhrLHZ4bOptWkTzomke
PcEQgtdXaftxnzCzxWl/NIzTW6Ze7ix0GkhTlBNfKUn2cFfJl/WxiowhW9j4C8LEhRWwTWb1P6Vy
HbVIsNO2/sDWTR7KFBZVLXs1U94/zpqkYm/Q0M1K3hSNgTTdewVtDvVC9YM4/B3ogPzoSe/mnhzg
I6FuoORqkihBZ0yYv5+JX6zgjUcQh3918ScsEyH7xrBAC6jJ9bDrFUZdhMc71eut0VfI0tQCv3rd
ayQEjVxmU0r6WuCymG5xJZwdcgbbClY1nQ1Y2ulmWFpTLWpli/Ctlh6sV9NQhhBcgrq1IZ1R6xk3
ddNLxTFb0rrBHg+/R7zCO80gcPtdDnj3CM9bLfQW9G6zZNZ7awIhAI5FNfj5DIHfOXKIfFXsz8ZR
yW5IJhtwSXaonjg3aoohJfXJTxtrJL5ZHlXkL2zw8FrxTgPpzj8ZTQ0GYw1HyQU3TwjEywqJut04
lVGsAPJZa5jsEG8tovcASEVgK5c5pGwDGceFYPEO09BCQ65WphikNvM9stWB6zdWXf7qrSXvFv7Q
zlFOpVDt/H2jqrMjNGL4vuT5VbHXsm8g9V1WrPkohTCWKlFN8Ek4k2QULxiAk/uyThN0qG2IwkxL
pPPjnyYV/+HyvCf/5gIpOROx9X5QqT2yb0Evs27wOVZTqkqReYR1NBTUnv9bhhmXT3fGW3vaFg3T
cdI/n9J8IrfWIRGRJK4gEmyu3nmBS77E044TFNkE5rqvrJGKutTEhqi7ZwC3Z6PfK+wZVDlpE7MM
2b1We+1W6uvXJswGmLaQeufUik9804ADNE0b8hgcz3Ss+fAnGsVd5xpSfuN62YYdDnY3eiObFXkd
su5vMdFCLomuSZUG4xeYQBNCP2ZNIZ80QTxZuXCavVmz7l28FXz2aTI8JjbSJWn4flKzkcQBJdtj
u3DSIMEH+l1a6hro7PFaisWryz1eeZV+jC3PjBHARA/yd0tOdhTeyfcdOrYgdGyPBMwUavQZrIrX
yXTQWLwi7CmafiIQtg3Ge7SOebJHrLzouqIQ/cfZuIM2KFVENbnM8hcVOMeqXy3Iu5wjuuazUpde
BAZvG71pLC1l+EdqUsoFYknRrd75cOupAfiMmlLOjwatoLEBGYv37ioX1RB7nEH3QaBaiJ1P887r
LG+L0o+7AkZzA2b60fdENJK/x7hsiTDEA4dIzjTLpew/6jlSzZ7EriMBZ08zozD0loNzmKFiP/S8
SEpHhWnA3EaFTecsvRGk7EAP9ietPOdyutPDzUGOPFDP9Fs7eIJ2fHT1UcMGTGMIkUdLDjEEjFfU
0UlUZyyTvDfwMnhANeIEhQapDXdBOgsSl5RRVjFyUb4anCl2jkY5NxYFwytkgbE3k4lgpBKysOKU
vtaZD8iw9uJ1p0kAaItYGLQ58MWZ8zb06t5J+Z36NwHvlba6ZBrIzk0j36oVax/lNvKH6borKpYz
vIgpkPzC5+Y2q80/hpiqQ9GbIZeFDznI5H9oeQE4M4uu/jeUF5wr+aECSq72pC3Kr/BtGbTc9NrK
xiAhxLuN8im8AXantrdFpggqf8y+7tj/Dmkd17pj2HBOnJ/Q5B6jsUYzhCChP3Bq1F2gnUSfPWjS
5OH5KOvDJ0+Ssfr7og2XS8at0CYvHQdCvLbWICqziQPWjGhC7KvTg9yoNyUdydZJKHfrrzZFFUsF
iyH5Stk1d1nZFpu6S9z1r8v56q/xyOXgcpQUxDB/wFpnMHhWQceDuixvOaCeaiugq0l3XKW5mD+B
IBE9A7Ue522gVOviPb8sY769CE94hzuRxV4BwQF8YdogY4Vlfjb0oQofW7PnEd5QxSfpbTa6Y4l1
uRnHo4r9vc84WTNhxP0RUegDnSa0UbTgqZLWkhEXjMn6iqaVFvKw2GRDF5eP6nHpfeRWf2Tyi//O
HwKDjr4W1GdI9c1l9Ow9/7h78NUC+CyqqPSsJbAY8XjvrvHF2oinDS/uZKi8x5Caq3EjDJQKDI8Q
bzZMgghmVQaeaoaUiAxZ5bXSa2Z9n3ajF+SHnwTW2SdVclcNd9+tBB6U+TEY2TZ/aZ0jTJANWLHZ
rX16Pf6knYDuzthiBcCCuhuLsBcHvZJbW6kjgF5WmEp8u3zNzPHz3L+fleU5jN8JLtfDlCjH7yii
PEz6tSEIo7oFaGvlDn4msCDaSECAaG4pnYy1+TiXDWpHcERyaTRSVfJOKnDf+vHr84CYRVT8lkKF
Dyu82bL7e4ykbRYtxM5F/dMtXjxrQIf8tQujthlpLXByXp6iFH4qRlGMw46uyTfFwesOT5M7tKtv
Yl1xfn+oD6+8QXBnPGGGEx2k/8rQK3yhsrTr5hQcPRsBBk1QkrMOBPGoTNC5/XseVna39qCaRDp7
rO6aDGcd7tKcMYHfg574CEx09jbHpYtDE3CVu0FZDeouQLWtdvUCpHOaMji/am0fNcFf9XWQ7nAC
sQAz4yLKVSwesHEgg4KP6XgGm4LfwSXsA2FXsU4KFKPBjWY+DCR+xUqUAU5W1g3rLxGzNUHt3s1B
+tEh/tLVZUl54xNd50wFtMJFDmXs5PQ4ZPug3vl32CWI8sdpbSzpsFUcRgdTJy5epWMee4eyQkno
74XNSKrda15Fsn39xXyPwpRQMCuddT+lOMQnB5Bvku/u5hpuhRBqfk6AcbxB13woKwL+F29UIC+K
pXaja/ibJ2H1rNDH7QwaqtCkupvpuIDKW02vvNM5VsFtZ0iLjR+MjSsPmndJT4JA+NB2j/AdI4vQ
GHsG2cqXftGifdKkqcUhtesz9CYtImhnxh1dCjL+MEW20KBslC6wEPavLi4Y1wksqgMlLrB4C1fy
Lwq59ZE8s60dhaZwOD4IgkQEwW69YNNDnzXy4+oOIxgRj3Zr/QjjigATAei1SuVu7JGmmn7Q0ZnR
i/E2IQqygMD8bWvgrIiDyOiGzX7eNw/2Edo0lLcmCC4qLDNShDyxlEIbZFGTlvZYgwIu+88is90l
a1ksKqYQqFdcvLC8PpnyOH0NTrsFwbpPDpKCAyiKNqcEXK1ifvKWbbmlDI2APb8lACzpMdszs45+
+qU1K8xCrRHhYWh0lzlLVNDrlSB6hhrrThvAlVhFTulPi+YAyZhHTEU6p1Eow2vsGTTUDrbBl33O
qzH0kQ8FCqPMtLFET8h0qm8Nxx5fwl9eeKZK/Q6m7nUJDMwvcdUgnHijGNOOhoLdaChTnSPy3VEy
KyGWJ1PGi/GTmAqqmqQy9rqGr5EuWU7hzpno2hJHm0LUrV/NhV7UOJ0obDxE2/ysASjL6XUqCHfp
NKIQb9nyp3pojvL/+5M0nDxXzmiJafz7ni1Wqb5PeZ1O0bV0umJtgnIAMOikGSD9mjxmDNGd1C3K
enm8reCBkf8WU/p/BpXZqLszp7WjtUwiFdt8NWUMQQGz7CwQsNaSEJw11g2M1Sb80yGo+v/R7dAx
kaQ+p+skIYf77sPVEoD8yq2XeGYfCJEn1Lu/HC9B7Fwrh0iJqvI+5giCtLqTWdHGCKwYcfvT1Dtm
uJLpxjdlf/yIInC5tjPgJv84yzHBUZ6CZ3pNnSi7UhWlOHvcSPrWe7VKaz3Zi3X/oTlB8OTJlcY1
1gji2VhkRjLsUF6QzC3C5drlj2qWIwOegftgRJMBwYDAr3UjB3Gn2ItnPSN+xlnA1huob0/dFp87
d9/HbxYyrgIPmdCZlKayfWJotVOlE8hDqROnlZBZLDxHbs+qdEne+NplsJrpTB3nGOoWIpB1ZNGu
9CuSIKFYQjxB940xUkZqE3n2VeOTDbO2c/p1sY5YW7W2hOSVv46Y3dcx3P8QXuSGK/GRNwiNG/Bm
OicpV3Q9oWph6ZUtCfOIix7S0groJryCdje5Jt3QZ6hqySkhssoeL1dNRshMHp6vXo+uK/emua0i
v9WLajn3F4vXFurLtkJ+b1CAMVV2Tk90gfH1illuBqC/iStbxfQmLqx75RRQcbzH9MTDVV3VxTlp
RwbSshb0dJYPphCgJlL0Zzuoq0u1zvIrHaaTn59qV3h1g5iW/mWm+lAzIVZ4z9Zl3Ed9OYUQH5oP
kSbdwUCKUGtAHn2on1BDST0br28W8rf73lbrxe4PXAdc+2zDhO/+8v6R3bigWnvCXRf1eTT6j3SR
svgv8Hq2PGce/6MsYqZbdjr6IAsNnkCbIn4BDSnOstVYTTV5XQc46WpScsr3HuYQS7kC1igKQxNj
qotXL1L1ZrkPb5qM37J65S90/Kow+rxy1P70TEDJJhk0xqQJekdE2CsJ/+p4nj8QV9fe6GKc3w9B
Q7HDa8EkvahqGbL6kIG0sDUchnC3wBHaCXhh2wLKYoC0E+YOq2+BujGzHobtMvmRjff+PaqYHIin
7OUmaiPvjhFBhKp9lOuc5xh3Fk2uNBK9hiuwKoBOwKpaUE3DyLi9av/XjQZ+1GpBfdhV3/ZmKLBO
i17swCQb2QXld0MJcJkTldRtaZvsTkx2P1/6xz9QC60lT7gZ2bEFcMixkEkEkCUHuE2ggGoFYX0E
FYqVWbTjSUGDPnEHMEf7aLd4pV8LdR2jW4p8+vN0WOh14E1zneFHL6DpR7wYS5SoPADo+5lxpQK8
A5IElr3xweWLnm2FyqTp48fX9xvRSbsTFR4xe4MxO+XQyFFzXay7LtlAo285hPPQ7uOME0tTY55l
vriX9xiTe+cz1S6JftcJGFKWFruLwnvZYrbmS+7Tjnmi5KYSjecnezI37MQX/GbmFLN4o62+Xd8P
yF6tM+cZND/TA0nY9L6p4/PnFGKa/Y4mD9FYr4lMdszTF5QtWDGq1yqLKw6eZXzugxBFhFcLihU3
NIoqy8boCIGC3NI11+36UByWYmY4uM7zuNUCiM59/BxHUwH402My7vtIqmAs5FmD+CyMouqTDldq
Cl4LCIBcHjgEE6Dw0GStPnmbXT+QWUIYDWC+yklE8b2rOB6/lJZDz4m4r1NvDt11VK9zfhkwyLuw
HL3LFaF1isf1EbwVm9VioffAvcxlxOPHm2QS2eaMLzpkRDg2CXv0lyHARiwupfw8CgTNsQuMcaPD
7IjXATpncPZtuc20BTcfgn7iTkGjXQ7bFXxRNp5Jr8NxaHlm+lN10ddoxR5klGWfRA/DQxnVPCqT
VwHRNL2gelcKFUwpf63f4H8k8/u/fnWMxylCnhQGdtAFwfHfxY48LVjsOs6chsS/fqUdTYaRUcpM
fJyYoZPHxJXIgtwYKsAthS0M8IlcXRjwvoie203T9pHWZWGJmfJfg55mLyPq9+j2x/64eepAWSMm
/dHv1Mc6GEzU5DBnlZMusYptiSitWfBx4KYSVg+e3k9EUAVTH3R3m425h7Lb+swi9rx6EDYrUILf
eA4NzYchEfDl2w7UZG6Cpq47JIV6TpLQW8Gd2qeCZXurBxXjbifNcx2cetQybX9QhuGGTW5PouW0
CpsBu0qLcTMk590c1oD1xFiJfacwLoeTnSAPecQrjqK4Rcma5fFHLZdtIZQIE+9+0FOK8FuKzle+
w7hCL/NgTcyoN7JJVFqfbFZKEy/Q7s0iey5bIbB7hLJ+EKzR7rk45SaMOHdBzP2L3eNWmlZpAlV+
p8R2ab4DdwESzrFnjYmk/kQ1bFpm+T7P1/slqdWDItC1+JXwIvdrglfS0etP75ViH3FH83od18Vc
vKve6IGUi6ra3fgTy8rdOBKXZAhBNkkZlWl2GjmdsF0gHqW7hfkOkI2QGd9iHrRnGf5WJnCqkyIN
HuGDq293Lb3OGWkGfZVhlEyNeo29NxqAjYUqUHhTt8yUbfOCRzKM9qZITtPHLm8JSLYEDVV5KVcl
xz6Dt/B8z6+f68Ktg0900zTq9AYDvQMjMotM/8qq30L/vvWJb04+TF/Leg7PBCSXHZKikj20U2E6
wYSeabfppjIlOJJZxsYw42YU+cMNhG8suqYaU6yRclPlvcvvFTVNbQ7MPYfTnER50HdTwY/YEtl6
+BdPZDFxtEQb1O0p2c/4r6tWM26ajkmYT9KrA5xlAcrhYicHpQjNefQoGSqepC7d4Idl6WyV2b+u
NZvzFIdHUAGyH8W6bhkvfO3h/haH4JsdFjrijQSCsvF5/yxPQOicHxuzwtcwkAOthESsUrJl5YP7
ELxbqKltjuziKwhPYVHWjIl9k+QMr99Bt/N/7iSjZ9axOSHzUO/FduHyFCvYueVi7gfPu+6e6gEk
rwgtGPUHnyzQU0e/RrmTUJOYcO/gbr5C+g5x8A1tUu5fvMjrREIMuwQrL6tlZ12zY8lT6rn3+AU+
eqEom54F3dUedtKAEIMM2FFFcMLAcOJudcPadTZj/764OXf3NKN/o7LjurHLPffgFqyAHwoKgszV
xlE/cgozb2cPcplYobOj7BlVWeQsjD1LRh5XD8lOS9v5lyLrJzFXd4H1EILzs+zGctv8ZsX8oyZp
6+pQqYd/P1ZQIlYlHP82hPaQIBeLtaYjuBpOjsVCsz7YTaE9en87rXiANNXY4QuPRU4WOybaD4ba
9CmmntB7XwSFjRyEUFmWD7KBGtGDbItAAwJ90lWnwRG68b22bYheG34UjBqgJ2nLMJVuyVJ6H67q
j2kp1sy5+s3RID1QTUuaHi1SqNHwgEG1hX3KXkY6/SVdSVblUbEQnl+laIdcSuweRJFGYV7TeRci
v9xaIq/LMTZoBfr5dMxu9JmaBShHASEYLWFpGnspnW+3Gtbgu8NFb0EslcfUA78PXiyFUVG7LWSJ
sdC5lmnQDtVwFZmdgyiW+JpOLW3bdw9l19lS7fIKxXg4Lr4hNR9aqTbnyGnBL0kmqXATKhzCp0LX
BEMd5EZsA3Wfn+iCQnrZvr8G8VW7y0CGywGPg8ehj5fKtvXChItVCL61OHngqeO6dDDNbOiAxgh+
MQylxySRm2bPa72CtZRxNAC5lslwSxkfUeDAMAhHIMuBqbO1XDeGgzhw8nsCOZNDpzUVObjay1Wb
za7plf/cWjOku74HYEvTKyNf4Qw9joFatwqD4Lx0+2WlgfyeY6Q/BBgO/ZHZa63OCbMOSGTpCkaW
NVH/K6ncRatAeVJwYKPghD+u+aJhnG4EMc0uZQzgx5+ujGn05XeedADEpgH7MTc0kQrimziahniN
qRAJV7JVnIISlHXKaC31GUabTyUCd0XCUvs6Ng9QQmVHH2Y4qt3rYM98tpsL5BTtHapJfCrEs0tO
aEkUDvDplkmLGwXIwqQ7dcAJmxyexNjPXZ6bI3ydDaK1yOE+Clh5wTdz1EdP8zjU0nhBBBA2d+Ie
KeBie60zf5OBvBTUTe/Qu5gjgF60kZ+0NhGzLd8TyXt0x6gS9D+VRNe0uPNx/k/h86Th5WbmDo6w
dEjfpdP+J1V4WwmI1HhcF1pqlrpUY2CAhOh39mdLueKpv8sXlENYXZxaTSwuhAfUdx8ZA/86LZA/
/xPBMjN9o0rZ1QEWeei8cYxCmYz32vIkHgtasC3LJKN5tBCaPrkaQJUjIiyJIiTiaCPhfoJ5vZ2g
y1yoriYuc6oR7zOMivnzMTenkf+iKgVSJZXRd4pzSOTnRaTYM8+Bg0LU9qCl78HemTfmJJqN8eVy
x0RiOXZVfvuI/Ok915Tk9JwpTGWG0MxrfH3XW9BugSABBMZrFrgNSrAf8VLAZT+Wa1OpLPvNXjSJ
tA90xatFJMU0nVwEyudXz1BdvKWj8K6ToEPYyBkAhJ8nFPVxjxgRQenYxyDBdEbSHMjKZTwzYgjT
ql1cDlBJm8AV2JDvu3wmhgn9zq+RnBcba0wgToCa2ZqimYygAQwua5xflpDMg3sNb2VDkSsZ1fNb
Ui/7uclUhTVHgdxs1y3DIqgxxTQuvFbeGB0xyZWuio7Yq87bBqd1j3GpeM1FjnW8r1rEQtI5cPdu
Hdnjbz2u7S9CKK2eh5sVOunILiodX+P1aG2y41wjGy74w5x3BSTVvuZkMnvfB+rZ5TUkK2sd1b5o
aNzqD4S3xsPFE0VhIG1r40n+wqC8+bFJg6MwAgBsAds5j0W2psg+ZAw4dTb8G9JbFwUtQ+2CNWeF
u/60kQsAGAOcXXFA0y3a02k8StEVuJqGxg2vJ3UUG0Jd7TaGGneN65yA/KglptqpPeUjfmmYFTh/
bxQ8x0uu+L7IKhIYj+qkfykP2+51sWPD/6Qsa2LFdDKmAW/F5AoArX4ZQsZY1f2K42Azs8DjeguU
CvJsOCFlHGpQLuIZTZrB6Kdtbm75jAB27RFGuD0h/94Eq+XiuFMSulR1UtQRIFP/Jka2sAcVDFIe
YXGz3cP4s3BHadZMZyI6fcd5OFqvXyeEDrfWgtHW5nByKK2QyjpnzId/8QGzQb8wrJdB1EzkpcRk
gMBxFUG6kCHUW92kbnDagwPNiJHZdzO4XVQdin6Npti3jGXn708ndmKrbrwwNoXk0YBekKEYe6zM
yY6pklki/haUjGA6oD9crkLXHOvQV1UXlGKik9FSiHxu31Y8K+Yi4ecBC2QyQK886JX9E/PXEJji
5H3184FfFHuP/dCV2bSblHmKSmeZjgnIQBO75pnmjxIM4AUDzwH/JzpVfdjqBpTWrNQ7juDPUQF0
I4+a3pPyzNHzyo8IgEPgMMJaRHuQre78KENzh0IPt3RyQ7KMNt4I5p1Eh3t+IDAlIIrvxctzuO2Z
38P5Lb1EpmDqGBz5AMH2iQEKeMPOZf6ewr+nPU+/33GZHD7XAhQzxe969ZwQnkQTd0DdGdk1+n8k
JNm2XpsFZJer1clqoVqmDuZ9DWUw80WtFyqN3sNMY+nc97fOUSkIJ6QRkS101PVbKgbOLv0lzSSc
MwXzXDbGfoXinJiL76+Om1bqT9p0ORbsLCHYRVl5QBRsWlfKuNw+7G2uNljXAKVLcfKzHpMrGrdx
5JyPO7wHcdQ2jQyI77FrgjCP0c2/9RXukxnRJMdd8f3qzGrHs1iuyQfy8IYFRt0c2WUAURu8ZlQv
6Y1+q0vTbnqE/3ZrB0QMTd4TXb4kOm77RCK9qGXTs2GFFJz2JkM9uXCt4A9CEx0FBq1Lk/e296/l
t129XEzdmvugDPLc81UMJ2cFnPYxVBswS6zR0RlmvDyPVTuYm6NfLclF5r8ZefjWWnyQFmmuH2Xv
3ESrmo0CUiGziK6H1aWiZcHTDTMZLDNfo3mzKS1v/Gj3urldaLGWIGD6LMPY7UEbVSOp4jC+MhmZ
8B6nK/CehE3MQegIo6z+UUT/+U8PIJf/N268NeR/cCNgTH9OidrteyKfRLgqzPXP9Zzt3muXcMuj
J8y2OaOmYOmjD1t8pO6U+5lzP9IYThnE8UVwwu8r9kjH11uZpNt2woazkTf3B604Bu47a9qyVVDe
gIPzpnIV3JA8y2xVFCgM69npdyT8ngUO2N1BuUQt5BstQzNGK94cdSQ/ljALjI78AH7XGYmLQGwI
8edRYFwHS8iZWu5ep4Me7Viw6ZpY7YATk3MXjdT/vf8jOu7tnF4kDiTITK8itJysw6THhEApUa9k
1sEj+TKXnDyiKekR1kuqFqF5BXsD1mkb6nkvHDw3fNYa/DvDQrgx9coZpIeQiCsm0r05tZLzKzUO
pNWFvlX/NWMX+QAWh1VYqO0zy+YA2ioG6iFUk3eop6OuAJOj1OriWlxb50YmG1A1eW+1XfCtJ1Cr
ZFRUgqJGy5xBGZaV/qDwqilJ+Y9zs88t/QmAMWFSMBQEyIrpfv5YNwhypfyndS6OHrQhDxgz3ckm
9fOyshdnqoAOwBHaxXSRYb1G3aSWTjXn7itB4lvQWf77XpyC9H5UmgEUyg/fvRzHj8t4RkC+ZHvi
x/cNpIAs6uDHQktx11ABeHfT9YMmsTvuwVOJmAXhOz1XbkcUqsAHFxudNUIm7t+yUCUUWrIQNQaV
y/LKZmj+W8jxNqUeTxpV/0i+qllCV6lGZ18CUlA5B58uyOtC1yAjHQcc6rkVysHaBCBNoAx4tCaA
QEyffPXI/2zhYVdHYeVaLTGgMUIKVmUiHcJnrGTuqeojqILz5lEmE4piYYetbNZClsyIMYJpM/Q6
hFgAsqe1NlrI3yk9SDe9VM5gThZAJQw7+uCNgX+hPeTLXt/gD0Z2XSxiZc3E05lTeX7DUepacl6K
uLLGuNlwQgyNSBDVrBhT1BBebHFcgoH/c6gCzAMbaQ2mkXiU4RTQ51hJrMsCVNl5WNGqW3H5XJiO
tDJ9Mt9jeDpcDcu4cfC7YuU6YrrMQKOuRYfcPEL+RbY8FY/Oa/TTThtOumSQAwAuaIRyasq6+9eq
34TrAGIQHhWnkkyj9rsLgZsMzQepjxEv8E8UofVWj9ei/r/MKKd3f65li6fFXWCVYD1SK4xkAhVA
kpCke9pNj7NPz5XDADnioZ969LOX3YncnbmVsQNgIBINVPfCyZMLh9F2rMwiywlWbfNTolEBea6G
mNl/+78buMJ2Rwf1SxtOfyAbOwZdjUB4+Qwn1fFPY1jNItrz2rV1UFLQnzFo/BLRwzNqaHDi7ypK
y11jK2wFxBSG0PyTLE1GvpUJBMkg0/9LUH4XgERr8elMu2pnjBBfdMQ9nQL+FZSMquZzh9DReKn4
jc8VV1ersyrVShpK+93dUkr+2w4j3h3j0YZmiFR0xonfwGm3AftvVC2Z0YgY23ZBHS92pBGR8ASa
SJJHTSATA8rcACI9/+3dnQz+HsiQW5vYbKIXxKeecLwhqCsVSMSWU7+gfv+dHMCmkUTNZdDKurEl
ORDS2dcno+NNT4+xiT+s4D1+p7Kq9m3QDwhyphudeRhTuZ/5fEEywy4uN5Jlln8FaUgxBmgFh7XH
aYAgpCANSvvjj1CBf25Xl/6Stj6nGSHOioEMcZvFOoTNB4vXQ5+bg+rsbVV5VVAqELZrsBC3fknu
E490Hczb2rIT6BxNKb/fRYg6XYgtkpWXFcsDA+d144gSxQ4qT0WORw8S1Xq4isoAIh4xQxIcxxKx
5+3Ymr52kgHdOAPw4OHnTTAEVstjR13mU3mPpMNo0tLjDM+a7ZnvS2w8GxOdMcJ75jKwd7xt9Sbz
qABjNMQGgQTZ+9qit028nD+Yh8H/4nWmG52FSoFMq/dV4Yky0hSUHX2+ssuMayzLU+5zTZyM+ruM
Le4oK9/cI/MHjKaYoqxXBAyR5mMm5RAwDQOaB1mQrns11fbTaleFyWEsvKZseepVqMGFfjQ+l127
FDsaUDkxsWTaHJBm6FSsa7CVTeElioEESo++aQkbgI+3P8Bh6V5G8wy4kONj8FbBdpc3yCnjCOPa
c0aNzVKsG3t975cwGw/bCXlzTQqh117eHS+aKCsHE5reNuqTRYosHPAGAWH1lgsnJKsd0gROy5zV
2iBQI4OKTonWx96R9fDsw/Y3s3SUqzc6puTbsiyN6zYU32j60/O5OPRIeOEDLd5TevUMg909zEDX
Cg7SDcUBl6EyxlWFVB2D95iLgDIcNOJ+Knw0oYlpr710aAPj56SOpHamrBNCDmjO/CoerGUlZnpN
b0Muc2HyICae66Xx0+6RGdg4z4qyw7odV9ZEoiEA27F5zFxiTPwt9nlGrwbAOO4Nm6KVCv8UNqs4
09l/9zFAJC11kGTLCKlmDIevDQjSrj4HLz2aBOgRo1bBEVtVUH50mZN3o9CR2rrtPiC9xeQuPGZB
WDCkCtd58kzFKJv6AHinE2d66EV50t30gYFLKGphS9eBVH/3ivWlgNcLX6AsZGduDPsfwMA7xAeD
tg6feZe4OZw+njjj66DneqzKtIohwS975v8DtvvFBxnfOsJ4x1+8IVV5GEs/AQux8EUSmNxxkOiZ
s2xb0jYodUp2qbPNWVAHxo8WqFonayf1u+dtd8YSD+9Lxu6G1tKq2gfGU2Ua4OZA9rKioXQKmT8m
ihoRKbOMFjgRyU1N4xa0U7yrqYUVESbmYmLHD4nJfo1MzRJbx0S7YoaL8wb8Yd3rnP7VtV8qoHOG
KbDtWRtqaBQCeCRlng/YAr1sds00JJ8bCeR1FlIrRlnLAp5Rl+0omMezfWrEHFMlf/60EkWwpTv6
jErGAul01BgetH5Hbh0fj/C70L5hI9oF8xsQ74txgTQ0af90BP6RRw+WRuqpPmARJh3f1xXR/ZQz
AV2SRVIXTMGYT124cE92W/mUWosbGcg=
`pragma protect end_protected

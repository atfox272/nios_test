// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ynkRNx9CFmFfjTvsWTFdVw28W3x8G0GrHnJA5BrvYoyXO5b6dnDRAe1CyBhZTg/m/vSpGRgRe2Ti
OlJRqEOC/PtcerEd9OgnYsZER/6nvgEVd6hrfO0Lr2uNRQ8i59fodIA2+JX5mdXCIKJ/EeWFsmSt
/jONX6d3LGMMv/mqocnVSyy2T+jXBappF2U6VQXaEWwWJONu7t4bBmC4J1SfB4Lpb6vLNWBcdgse
Drr5VUn6lbw/sDBn/bPyeKXPds32391sfMusFbQBVZOEzZP3qExMq0bjUNEMQe+E9W2kh5eOr+DC
UT/RmN6b6K7mQxGPfjmk5HEQN098Znqgkbi+kQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 12912)
CpZAsjTDAyaV85yRP5whQDdV+ZjukRUbkiqkpH/Hw9FWG8f1IlHHvkBeYP8F5lGDww1ErOX7JOWy
5zrJ6EtVcji6bP8KIMP+wdogKdUtClndYpXjQUly2bYxjsTQCy7fqIYSGXgjD7vU6B4O0O7CGb52
SftgHJCF1dp9REJxNadaFLGCqOLqf4LgR7cNN1EYqziYDQllN8bdfenbDTfGY8pmkYKojRK20iTq
64///MR4jIMPQC+DiuxmEUB84hzjBhQF5t+oAjIQMvSQ6dA/Rs1/HZx72Aw8DlEH2PsFRRvrFmmQ
fNMl8MnTh2Op5wiLWxOECGr5MTf+n2z+o+P5h3oJawgiE6HTcr+iFIAwgNxQqXiPnNbKsHDocMp/
4Mf09P0I5SSemUS/vUKErA50OhEuJyvBUnC8XBmkZtmlgHJs2LfBztCRCYkg5iR857Ek6rlaaNUu
K63e9qDqFCZUygOjoSe7BVsgeg/VTyNbiTQLOy2hf+NkC9X3RQASM126sTrKB/flBsDkzkQNKJem
QERCpo95QK9vP9HMgD9oX4bVv2U980AjwvdANgf6hLNoXMyaZPczHfYvQlA88ocvChPYwulnRzan
lTWRWf4O2ujaB+X9iJRSbLwHjEu++ZNhtJryoypqN6Y4/hPti6xGLtX0w/sHJckV+ZVNzucDM0UM
l9hCzD806q+S6X9PtugvtgrSnp09D8ARF75h6lPwOHdOkBl8WE18cdk8jsAFDjKkhS5zTn+OuIDe
s/kaDzCcuHZGwvBTpJoaOmv6iVPT2rt2Q89BHeoFK7ICTF60Dk7lIqv00J06h5TjRccvjfQ4Kcyp
djz4wZOlumqJ5FRLDaMOl4KI1CaiT0O06ZX2Bd2Pj2bIIZgJeuu5LvzhxB4+rwgOznGaEHiv7E52
LR+dWG+fc7ZCZJw+jYx3kMAoh5eVDRgSIYvnhS2DhuWzI6J9hKT1n1jKJpMZtSgIDR3qz6ddyR7/
92EOOybaA+FBLT864vWcPDjumrmDamA+RmZU/KAQPpqZaWnu1ES8EK4ogzaTIzuXS2a4Y2v0nAw3
B9pHAHIeFSz6KgpFTw1+tA6/NUui3pFZQ/B8blu3alyaH2Tt7v8Nwe+M+3K406PM+wXgDBwJKGqu
zvp0xBbclL+418roElam6P5snncD5LC03tWrFbnDzFjZkPSUMXbe5KmE0KL6VyV6xvuANU8fOrt/
cAc0Fplpkb13ou6PN1wj1636yseHcwNX1E1VZYvLZWl2nE/3E+K9zl9d9MFzG1aWjigzfF0z2bGy
YOcuaFbMgCgOJdXyMHV2xPb4qEWRtgZvY1EC2/aetRhzSf/u4b27PWoPggY2d2SNxbE/PStqrFrH
+T6f/5nj3oD34Z0aOu1TYPUmgOh8D5uMb0xrRuPp4XjEUWpl8RoFrSpHGRb3T8KfUpEzt4kRQ4Zl
OuCmIx0VeOgX9BtctmtTAAZnH8tJyoBAhiYv26MOFmMgXYv1vgCy01cMdR34R+pd0T0xWpB3YAIk
+rQck8MQTTtYzlfkG5RQo+7LJjbK/OWiQVAbjSXF7PQu7qV4qWz9pFWA7XGAT4GRGMmI6QfMNbGn
0BqbdFWBX3kreJoVyEQ1d/EbhFl8b0hmUu/ycUukOYM19WtYTwUDCt5Em6SJ5O/WzPOZfo00rHQc
MwU20UVlYZG0nTvNAzBWpz3JWeJTEeIldu5bpnVUlxq4P11E4s3ODGUoNlk6eJwFZueZyBLgsVz1
6CF1PUq5R3MSIbAUCyr//rOHZZpCOqAeOkRoIUVG1Mh+vbwKXYS0xFr/eZr3BtCSawlwEIYnaG8G
Rn/IVI3myHvZR2fGBdt1qT9cuUaJ2M/dtZrGrje8+rGXnHBZ7dTkaXPts4tX7LeSZz/8fwQ8/BYi
On4cZRQXlD02clDi8a6OjR5Q+Pv6is30T+CYxZqHfIvEEQbIXpvEZ3MlHZIiig91QkzRQnniAwp/
+Q8OQuE9YY0aa1oFaPaNxSNQ9s0F18wXIPdtdToq8yc7JgGrP9QTe3JZamAAOMxO3XvhxsmBfXEC
WY/+eqwYiHSZXmy6olnO5/wDEFLLs2eIXcZ4nvTddmYxi1++WLuioLIFMi637K+P6EnLT4m+VjAR
UxrTG+PnKuQvLZsd8Xl5BZ7Sw2d4UGDKJTKjY6v0fyDwq3U9FDuSf+9oA5LdTaXDiORSw99NewJU
LLKXyAtxe/dglPHz6fyCxUwVGAl6XAm30IFf4+JS6R8wFDeePQ1ZcJThdbHJXXv66TSFUO3mqqEV
4dfpZ4HOAWG9VvZ0sWFKHXoV7eIx/ggFsH7/6fAbydlkB9/QFVvAEWIzwJRvUyk3p9i+OOX2yyCE
EqyMgIF1hJnIgg7Do+sV2ZmKRSkqjm7mPZCYC98jsWILmVwBjhvAfrpS3vFl+xqPez8PF5U+l79Q
IKEHnodNTXX3isB4JzRemozA47oj3vNw5EFX8G/mkdhX5b99zrUjqPMjYecfPsG0Nm/knZbp18Vv
WEbJpz5yAvSrqXV8avkb3tjGcANNp6USEPeFcr8vQp1Zx+moJh1ELZWZiCAMXbtpSV22dT4F5YjV
Ev7S75slTuxFCSZLjuDn3yq+wgq+x5eEhDl9INZ3Up8Jdje4QVIvx+B74HFjP/tysW3oqD6Zsvnz
jp4Br26X2GgWMMnJn2EfbdBQcRzSiYSSDTYOj0Awe/WtRGHft4MA7O4tMuMKDGu/UCXPUMYLAH3X
OePJk69UySar0oRES1M8oha/nz0zQDVorl9v3HFPFeK6kDeQ+Z/S5IOvkCfkD8qmeFedulkEQSEf
0DC/CfoLNLNO6x/m0ENuk1a8uzSmScdgrShnArMZKOYRKn4HH/SjjKmogCmgjsfTRET9LxVI+unW
NiyQWOoQLmQSTEX0leX+KLHxJFFZ0tqDnJkt05NcXLRBBcLJTEIu46CBQKrw1mQebxGxA94C51cg
4a2tmRIyxtGg1sY+2I3aZJSdUEqY0K0TPz87s1x2LDM7gN+ei4yalIfCZlMEWL7Ae7zyZXRScBKO
HQl5tJvBLckZn2VqNZ0tQa2+36zeQCrMlhBe9lGd/aykoInBhf8fiq1N2/LJx5yt50HbjiBLMJ/g
Vwn50YoWMR00J491MUYjJOPp1XF8NCPSzHUyG+FYrDWxvo2D40QV+bIRQnXPSqbuVIwXl3jLUidH
RXaXMwcnipVny14ALOBseI+aqF/jbI94kN7+LxUrQHgfaYDbu/PelMaGwWScJbTET4xlqEeDdq+4
mKD3o2gEXTFzkRMXBOFZv31rprX0aJQpmKf1D7sqSqCV0KUwbXDS2lbCJCFiTvkU6NxPxVwxdV1c
1YPMmehWDIZN8YkLh22Hwxycju7VWjT/SA7QgPLLn9kN8qc30TZDE+JEhd0IauhYhYuNbLHih14G
CrfKn/bDVPUkrgDNI6E7MODTU0cwqVRb2DGqisvjTqVTYTf48WMQ44isdKv+ej6GsWyLpseMLHrs
+Ent394T24dQ5IYzEeGSib40ffafoZzOAlKjycgkfXemQ+H28y+AJS3mfSOImsPg41lIR6PZp6V0
U0WOpASkgpHZ3RHmeSswcn5FOMwxIe2Or6R1DCSTG5y0wlWVtnzYBp38LPP4fKy3QkNlH/GmAoTh
gwv1VmPbwK/dZSeaWGjeRaNtyM3f9HOQKZW+Wnu8xRdJbPW8vbQdhmEJHviYYgXvF7tzmeMEF2rV
/bnVE5ZHhQsfCqF3AwOrBCESRKj7lPKjuXCcG7CuyZ6EmzXA9+dYUxdEdIh4O/aOLnVJS8P+5JPY
lQ0M6sx/MaohGNIP4c9xT6fHUF72Owy/pz0rMxM0pq0Oc016Ov7YqmWEQI/3m6GGnotS8B6sQmRl
gAtaL2me+YmQxMCwhTAXvUZj4JsskQQKSI47RgUf0pgsDJbglRX0Xo3BJmF1CFguy5pBl/cDPebD
So+qHZ/kN8+VSLUOr017yn8Q4GxJA84wTd0IsgR5054JuUMH0jAQ+LLDDDDZXXTPTeFKngInQnw8
1wxNjZtvKdMoiT6wkuupIEOa8b5dD3pLwbUjtUAQmHTHHS0KtFLhDXUXxLmt3T1cXq62rs+4B2nl
8GXkTvdRW/oxwfuBXzxjT/oLsYpES+Fkb7sUfAUNaOZfZ5bHSY2iGNxp0z0H8On4DdaOjRGsG5Hy
CRJfD7tA2BAl5raxVr1jkE/w35VO96VwqeXxKoEYHnuCF0dL2zyY16HItRKYSNNO37+5LuvNzsoj
LUz/ki9HlUD0meC6EuGxNn/fgvws9p+nr5D4xcTPtMl8iU2jm+DmJukEc4pZGtX8X8Co90/kWQ8y
pu+NDrW2E3JwA6Ov7Gj8DvYlu7opVZSWTMq9p5KzFo4nQbQij+JUqewpociwRp8a3/dWEVTzdV1v
6hBKCycJg61Mbf6MCqQ2wIjyg4miyjAmBNm1HoILOSN5Pm7h0VY3V+x/o6rRWGcn1v3vwN0XNgA+
vXjzDFuNLNogWTMaa+6hf81uRhe2QmwNPsyYFGEI9hBTk/YI4EeXSPTPmfUVmF4zbch8d9bSABeo
fv11peq9g4anyLIVmwQCs7KiPZtJMrrQUBTvaU7rfiFDZ9wXgB9S0ymu76DqcRTh0x700iIYj8Gt
HghCrvE1/wtQnTAOUYtowblJ6lPDiGUr1yLamYhglwc87tDPuV1dtRN3ESvJQcYyjSD+M9NKgFSV
kBhVCBh8hb3+TDqNdI58SRlkuUtyOriydVidey2HGpvE03Q5rne64gzKDaPeAIv4N9rNQh9hrToW
87BVx2eTYS2wWQxu+fXPDn/3g4ZL5II7HSNgN6UYG2RGpP2Et4Z0Gibo/xjwcX81J45TESmcHkKL
9/9ieJP3lHzS/JrO7r2jeYvtRWhhu3TzEQvL1PD6BUswJRNRlE4b2QwVuggagzsKPpaj8xNy7iwL
RA804kmdoeIDjskVsjYfkCJyN/6JZ/4I6FPvKETYwEUxWyhDhk5hrvA/af6eKoNnkzAa5pq/FRJp
Zm916j3t1vFTly3XGXXGPSbTLFtelZCIldZ/6RQUMkSlcB5EXKVPk2emhuo3QcgLXcnheeDMRuib
u3weGG5hk8Bo6gNLUyAyqN9GmoPIa3LcCHdKjAklVp0YKhT/SNzKCryvNNhDSSzQ2CoGWjsTd1Ri
IG5+Xyp9qlNiOUixg6JzCJJdlWequfL2w99BotwtRiLOnCc7fdInGnL6+CNV5rpeqYaSnRBr0VuJ
cYwEAyc7M833Xx8zmFifnwZ5V5J0IxjMUPuCnwtdFzKhNv4xaRJ8HUGBbNoNwDOTYyHJNldbUGcS
Rt8j4vftHw0NJmIRcAo89+McI3k0XcENDWQnBrhrmW5IE4prfaSx2L6S/q73NQdoXFR7Y30xYSqP
lfFBcXleaAseP3vqurisP7ANqYLrard+nd9yknJ4IUJqON06XeksfPL7PGf16SYE1mGBPngQkjXs
LfIAyvluazfHqtvF+hueYVQ6Lc8FTaeUGOHQQzRIdsA4zBrghLPxzqdWYj5v1eIrME07j8qqt1o8
PXT8RYoJ6UR1d0ybc9bDjCfVgQYZ37HN2vGTncnyFYdkei2TD7ySuH8P95W2T6rXrXZnAWHDZ3GX
W/WfJ0gGTw0M838XT3I8ay24ZKucuJLCz9VW/xZ6Rsl0FSrL5RdHg/ceC7FrFxBzbw8bnQK4HqLd
COQp+ZluTFSKEXKltwm7zwlc8Vq1y6E4tDtI3nXHYCtQGNZq4W/W6UnV8Mal0D0IiDu8tFpu9fbO
jnicx46xZNE034hA/8WE68reQm05pOV4LGO53N7Q4bzQPyR45VzQyffW6UCSC6kMfhrJqulCQqeq
s8v+tapBbMWVovzin9IzAjWknIx19opxhrkmWa/Lt0Fe11T7GB6vnPhUpq2EPLosmO3vPXGqPt8G
NWaEyWaUNboA6NKmTKTYTXUtv4Axyr0RjiGhKlwgAnA8YiylEXZvKSqwiqE/DrRDD2KIPlXQ2Q8F
3f9C0XdgOqveIPK7Q2QpntuWDxwFYqKuOs5x1lQGmj7NWKhQ8BzH1orqEEGn2IoymEilqkLvNzYH
aC9p5zHL1Qbv1k7gyc6QXKvuNJQhwBO/siHjuP/oHNHzWs3d+pPgjpuUo6bXYF2di3hJFZeHlVIh
gAM85xJq3RqO/NzZVqgHA6oNMg+QphNzXJCTM650GykU+EEXFfKb/lFR/0aTr1jFiU1A2Q/zWAGp
H1ooCdGJMgR7FpHOnubRS+np/w+2t5gJnOK5wNc9LRdBx3dbH0b2y+dK8fCPhENt6HOT5QINzioX
Pc0KLyIaWfTyU3QfX7DRw9oqCHFVspmm1xGyNMHLRw0byvAilF5fQktVpSCU/klJEUtybLT5N4aT
+H5BzFOxywW7qaGCPF5eMWR0eU1Nw3VO5jdsWtEk2oeOmUnb3HYMPb3koMXKbt1VOCxmBvfsDh4P
GY12bgL+YmuU1QVc6WSyZkqVjHUfFX6c4/oqk5DoQ6p9s0DuZYzqAP/k/LRMKfTQJFxKtc8BEK+X
Jo63q6k2DjICBDqrI0zYwGBNBh5gBaWqK7BEaulVymlIRX89X7dMjqhU+Bl15rcicWMo1S6JdMfc
r4Zg3l5MbxXjWh4eosS0I37nBegtq1rT8fOp9+Mom5Ri7PciM6GcFq5oD32V04rjwxlh/yTbqMeV
13oUJNycV2Taw2ZJXb989aldvDJuMwaMd9sYqpBOnMG/2dEkyLxiQqXw/PKCMYhMFRK/tC26CNVf
yCiej6EtqroWueOyKHq0ENrrn7KTJ6W5SDDD/jASpi2bEXqlVTDYzD6WYromNayVLp8sy35BdrZY
wl2/omeBNsn5/jk6ll1Z9cUmp8lOD8a7FMEZZQPmTVZylkGJgs1x9qkmlBfIzXNO3q2IjvcgYqm4
UiJYHMqU5KER19gZ4pp+RfOGtv6NMOyBYJ1FYx3l1UkKkb+3VI+9//zOMkGQwKBSIh6Efd3ntEJv
0qrqsjNkSORST3yLZ3bP9qvZ5QWbbD+XLIJ/y/SKa0rbnkcyYlCnCojU0oaBmwbaZTRuwPkTnzfV
AKSGjzu8bY2iVEk0rB5rx27r+lliWXQu0pAUyicFX6q3L7s0NTbvTw6dPyOEfknfy4snoywbbFHx
bkdzAHByxABLljh0pWLME1cxSTi7mQzEYGh4IyIM48/estLneZ8kMWq7IGW3MdyvXUoA3YZGm6S6
+Otdl19cmIkHTwKj4yM47w8awAIGD7RYXJoQbvRfTA4EttrnLqE+hq/Vq7nroQdeMtNqyT6MwUlp
SkC+jFOKyw4yidmcBh41upqKnP9JNt4ywaMyQpXFHmWCc4yfvSct+VbU0Nir831y8YehUK1Co1Jj
DjoqrVHMfJxv+0vD2YNThIHp7vv2Y19YjebR0br2LukHl5FdrZBhYrrzx448ptK8vb0ycInT/W6Q
M2oLXigwMXT4J0XYWcnC0RX7xkyIHHieUtPRyGsBUewit3pTObg9FiGmrzlTNohlg0Xa0d3b1I4C
+EEDSj71s9WYdMWoHCcC5Zl28R+QUeZ7l0OY3C48eMTVL+4OJlPBlsmtUDonaNREzsjfLCuCbvHs
wQebR9YeEAmF2D3adR5kbupjeqKxWer7x7s8EATZkuQdqDgFEB9I4EZL5fuf3XU4uaC6K7iHEhBc
7a16MRnwJqzqglyTF2bX/FkcbtG4wooIYkC1/gC3bCC1Q0+DeSPUDsvKiTMpADRhgcrSfdokNVfw
QKR+nrc7eTInBh0BVtLrie6h4MpyJvOxhQTjVQpsYv+vrseV4zmYTATnkx0TpYU/3NuVe78GMVuv
hj1BJJuJdrO6TR3X02NZ0kpVBwq5Phq1vCShear32sMOZqrz3PSwhG9zynCr3O22T1LaEfz5a7xh
9Myyn+UlLAptY6AqqrojVh8kRrQz5zQy87JRLdWGUmKyMsBkr7+XYByARPTnzI1Fcsop7PmEFCZ7
RMSY/HOucodeRGOnaLh3lHDR9n5iedLcwX8jiFmJnO70OxAdR40IZgbPl/hBv+obwRkcwMDvmOcR
22HxncE9F6OPwGakGH/LOh/241gDCAeR5wQTMtyYB1M1c9iRV1W58/A2g43Rd1ZQMGegcNnsRv74
fCm6jA160dFLpFu7klw77g/ADFe3FDHYrDhDt83O6CapAb0PfOfcyeNCebjdcsj0OZaq0WjYOYRb
uWm4dN2DHdxlN0dfnC4FFeg0fZw4oi9GkXhBSduiAQLMoUNAy18ePHiRdb22Yzl1FXh+kX1ipeJB
nQsAeEnjZgws8E/5EKFjPu2dxbrmrnH2kFepUH2GrQX9BfsNP5soeZxd/B2SBAv2K53JHlIXbsc5
ukl5f/fzQpVLClYQPH/XxSQKUN0w7poEysrQu1JN3gZ8DsquCJ78l4LQ86ltXb0XCBmvZsnvckli
dSxhBlCqv5/AGLGySWowU8gGI+0v3n5aRCXnkYH+crutnaZP94Fd4m/uoE4A3Uv2vxcqR1+I5oSe
lO34l/QQ4EbOjnchkCGM7oip9os52L5eYKeNziPMQNy0Qpcdm4/uzH9XfP4AbRGjfMrS4n9f9yb9
M8uajIz9VcHFygG9jLugbBuN8/Vb15WtId3hi/iby7Rp2onkKwJdj+Dz79HhhfCaTHuNHMeRNHzL
/37hDyS7chxWfCNjQW+/qXfTqR3R1ziPJ47YwNifiov+Z3w4hhhvzOkCYSuEczE2lWfXbn3zNIEZ
DunThdwKGarz++PzDopn/J6PPuZlI/av+Jn2FxGcQqTF5rlPQMe5GT69CJUrjZ8zz5mcGhBONlsm
84ukRuA9TGdX5TwLNTO5ptRYvgUePuyyWr1VVSJn0rZ+awybIw+gp08ZFirsXX9re6ykJvsQxTvY
TkYLtN+ZFSKgVPPWP2HLAXDKIaOrU+UrRFWFSUujFIT1Qhy55MwENxbuZAKTUX75iWzQOItqdjl4
jTfGiEkh5h0/5P0UMqFGUnw8Aqt/eVzIOz7zRz5JWSXpYTFXHsaCcyIhGjHhP0krdACZ6HgnXoLq
f+koSGDZ/ai4qFvVNrWTQuRPuTv/izP9qEpYCIXzqP7F1+1J9QCleVpYVQ2xL4kDdF6O+qmKO7mg
NnQETtqyp7kLS1LX3GFMnObztcd6mdM9lnvDRua9g1ynm3wCCBwpHi/z4XlUU5cqzqO0vSRZjRjg
bqN5SoP6gy5dFVHAWTcBBTT1ZAg7zlGvyZF97R2FbR86n1p/9DLUNOhJMHp4nXxp6EKwLM2V1PO5
acHenJSXQd4aocFCCgQUolKh7ZxK+qACOwb8wQ5iR1QhZZu595mHB7rds4amNE+UWxNPOTt971Yc
n2zbhSs8x9KC0tbp1XgHOx2NFFNSkEmLxP/XgrcaaE6/rFdKklF0RreqzrkJTLIiO1+D0kPFLv/x
LU1FCVY3C6rghEZiYIoTTZZ/Nsl3flJoLEbmBfmCu8VHiPckLkk6ashRwU8S1eznKIBFT/OszqrU
qdrcTTkkq9mAEj87eWe0y3qEUebAuRSuMS9WoR9gLi6FoVXHTlYtbPUgdu1zuQ/6VGHVGY5QpCS4
QX6L5/VN1eRuZbg2gp9f/6r9vf6kko5mpCUlflxV85zxMcM5Ur8oOFQZloYEp4CHFqf3lSD9mZ+h
jvdu9HsVPKx3EyBNtNJLBoPuIkXxL4rnek6b/nw4eIRdY/mg7ocp8pMevdBfnjW4hKrl3LgPG4za
dWJjLFYIl2+DOr2OyXtvoyhRGHe4Gxm+2lBCiI5MScQnvNw/tSEjdSQ1egsH59zskE/2tkJsg9o7
EZf3DlDolXXgDcyUX7d2nYoN7/pm7bwP8Nc54+s/nIyepE7m4xPGzz2f0DXc1Cn/Y2pHwvXzWE/n
JCce+pTVHINCGDkoGkpFWqV/KN/Jb/xttpmRC3Jy4nO9+mIEdvjRehp2bIVP/bfV0jFuf6GbaiqV
hDBSDS345qkC2YLtjfJJ5kK8UhJsi9x2+0PZhz+PViS5MlhnpzSkCa7uD/1RLDNe/8CXJdRfdk13
qChyoQcZKF88nKGqm63D4Kkqu4I9xUBcsYVl0OEBfaEhmusa+OcgCcimTf62HLHCVBB3OxMXhsZj
HalCBYyaIaJbv6s7lECUHlehyWEFAglTINyj7t4ojSedh48ppIDLJ+LtCdNpj618JT71+m0OZ9ac
tb0Q8KtXmcLEllFWrRrMdm9pBvKe5Jgc1+MfHJQgiEMvzgt+XfCUlo/Cn6xI3DQTeohsH4q1TLig
wlbHqi+nU68LV117ICanJhtanzADDesIR3c9uOYVaYeD77lO37AkU6lBMP7sf+S7iIdHOA/XWpmV
nZ5mqmoL7agsFgAayzgH1WY7hdHaPi+KiPPCF/Z8ThF78tq/CFb3nflq9iTBWSvYKH8006FOSbKe
TnsIiG/e1FaNjq+gvmMdw85aKUM0u/BbrLLcyZfeTLRk90RolHrOR47Ah8Y/SOiiGBnJHV1Myf/I
fh7LElnYuA8lFBtT+moyFTJf5yplyza0yOKi9jsfNnUsqenOnmBXmixG9IBv1vH1b0xcLVP3RXsA
DyvgsBeSH7FKZaiAd8v0KOaX5uQesE5a5IBX4bgCxknFYLBvCv9ckpMMYO6FH1aHu0NkOjJLYOE6
BC5sskxJxBXB0HlNnbswCaJOZ57noSU6yMOly9J+k0/t1hv6GbakvlSLEsjADPZajikI/ZfSR57B
G9c21lcLyQ99LCETaBrsFIkq6/T9Lxr62WDZyWu0yyr4g4bRaiiysx0PjwwbVJrQdce3KqxTaaso
67lkD7cgsKtzDzPfXqTPHma7NG6klQn/3eYNzdoIcrEYyNa2UNn96nv6Ii79/eopuV4XBGMKFkTk
bk4HmeWFmOcWW4o27/MYSzBt4f9T9f8mFWnFrmeBOiQhsMnI/PMRpDG+Em4erycoBPnC5KK2O2Ko
TLymGCd37KZQ3s7w+eShM3Nn8rTew7zk87UMzINWsSHLknLnQSHuyU1y5nzYR/aIK1fdCwggamqT
ZzRswFikj1mxvGowH0P0BKVP/ZTOufPIj+gXLlnzNEeRWy7dxHmE0HAo+ENR6sEAJgBu6bsBfCiZ
hdMY+weCMuZDLzhZXnoCoTI5ymM8QV7cS2LMFMQZxDJXD+YBh5dclCvLl8VeHbutquzsFDA3JJDc
z6IV8E1aRv8ksEUZ77pCYMwJaYrlvF5QtNMOgP8p8/30MnpaOfvU1Lj1HeaOMk4E9nYEZpaPrkQx
hhQ+u2vR9qUzgmZnq/8ci26BLQpksZS8zE+DmMd8oHrRS1Y30ZiZSLSoVOGIzdDuGD7UfPseOScP
wN75TcBh2jY+cDGCZVbXhGUPQJTAa/Oj9ZAbuOVmPYnkHms0VmaQzSqhY/GXy45STUGX8/A5jdGq
vqhhBzdv/Ob5C/OAdHrTC3ZuD+zSe7Bm7HweunCTH5PfdRWoCFXs2E4qTDWrTBoS+pBS7V5DCwHY
KFnOYPJapSvzGy/L3Wy1BoMZOLQUi/oSIvvPLyuDbTLk0jjHo+RWEX5t76mHdwzYgKuoYtp/MmpN
i5QkMMNopkaFTUr437UzKsp9KtrIun8D3dyhaHTjUhJMEfmJJDKw/JbkRDxkYV0OmWBcCkDVGn4r
Uw8gRfzKOrqDR/LUefwZdKz95m94jbkizOqvwY2yrD3eS6x9+vaaErAxD9hujjvomCPaUG5JrFDV
E5pEw3xG4a3qsJECA952igfSKQ3OXdueZpPhAz+a3p2CEKXORFXrsPQRWvBka5U3SEN9j8vLOkUE
grg66nx+pyi1rRJOMQIVzwn6c1mCQH9oe2dlcrXlbJhQiCFgR8xN3vmmIxvOsn0+OIfLiRR0ZIkr
WsmKcs1oVXNXD0ro92Mjpg0aLgvRCEGansi9z74dQ4zdpH+5SOSxVpcWrepBBvINhdxNENEjzYko
/RF/Vk4AWk0Yq0nYuO4FlgYbIZbKgdhubCcSGARtBv4p4fsIRT4XeczEG8RtxrNHenbS3NAFGtRW
w//tMegqlOzHr10BTqVG0BbiTvAoNF/2j7Vllv2dk20pBG4jjth9+3oFjD3gsGmILAsZnJ98cOb6
NCiOOd8CpjHsnpCrAzR4wynHyoQCDBMdv/r8s0PDnPRFd4SczIrx6Ta3S4ZCVUmA0XlZtZJGXxnP
mA0inp5vsjc1SxQztUA15ATHHPovDAYbAMyU1Gm+JHSU3EheTDdyogFOkYsPs5COqxXTERW198dA
qnA2Z8pWEawAN+e5x9ZduVcgmw/kucM1jvOkyBpRO7elU7gIyBopVrj7/kFBSzcc174z0oohc52P
TzPlVyIHpOHpHQwWDf60Y9RulCy9rSpecWpupADNvGT9wH9EZBu6BHVFI/u4TzSOZ0CbVIfwRVbJ
6EaGBoPeBtFAga7t9WCUc7xbCWZ1bKg2hpLS4C2wjKqQtsDItJ/obZJIi+U3VracozQq78y+wg/E
Ld//ql0zDajcafFwhlPLe4jC1WcE/TOiUuBHyX4fAsKnlnRGTLdE71pkSLcycRnIbP9PeT5Wv8qv
pb8rYC0q/zJRLUkOHdfjADbU5hckFzfpNINdyTHZIeybYAi67TWdpYt9nT/vSi3IchLEq6Q3b9Ix
9wkfHTB+2Kt/EpQKmdSV65Ix4w2CSWN/f3J5b3GxBqZpj7zGg5lWDvHEizk9EqDo/HVhHtAa2Q9J
SILfX4IFRIMFi5edOSk25eZhB3rALR4u4b9OW+t2pqB3uMMqDwkMFGtr0ZB048i7sUmHYfw14qfl
yngB/hYT54iQhlm5Bh/hg55SzsAd5m7nzMk59sKAVAgrE9WnwZRRc/aCh08VL9eKFu1HVNiJOJTn
1v8Nd9gWPsEMtOEdOWqMNUvyd04G0SAz0WRi7wNCUcq2rBtWktP+J2CJVL0RANpcI8WzKvF+eo2S
cCoGvw8bYStDjZhRmTCjB9DOgOh4FFH9LPe6dnSKyNoDHL2oI2vGl6G9ewFOgmrko++P163lIRam
//Nm14uoYkKsdy8lJFY4qCOaDCt/FUUEfEQgRBo2oP3dxM0+FWxpqxfqBHsgB7G6SjqLxUF3dJEq
QGIzWdbLT8GqcRua3geisSxQ0cycoOZGrC7x3HgjqKS92OwWun4dW67K2VSJURd7c0cBuSKmRi4x
BKRWCQ77REJ9AEgQbYNicFaCVQvNmDS9MNC2WOzSWSDIGF/fMLft5pQwjoKvZwbRWGjQkgoZvBBE
ENSEJjRKOyF8wft+fbo5t1V0ssLWKMLCFwSUZZkfaPoeRWHDvmLsRvGz58TY9oMY25HGSX0eaPOx
UqEcW+gvb9rEUsMSeOXY0jzJ+uSVz9+WtBLbbJFsQiz+F8G+4zmgwbR4yZqO0lnHIzxceqaShC5J
LUp5ZDviKHxlgPuaug/z0/801vUkXIAwzDHUQUgKkFccd14CEU3/v7eQofJNcFq5R6Hcl3LgRuCE
nfExa2sqQZYyGD12VhF5TxCaSQv8ifeim8069/ERNboDq704qW97a3CVsSNWSiXStZpy3a61fMF9
ohZ0opjCmrcZ8h9d3rQAna0A3kKdtG1NE5aharPvJCcu7MpMk8aNzK2tIBx9w2mOSo4XOhClPUPo
m6NuM22hJKjHmwM149mbxtiLHbrbAOtr43gT3U4bDyEiYMr7Fg/KBPQDEUfGIbvYSSt1JlP1mJna
+wWkR9FAbgvUtpMD4W7jwXd6Ih6St9Xh3yKGCki8zeg1LWE/bs9ozAZSemyMmG4BewaSbZIISr+5
e1MROmFqy4Apda8pHZCm2x8twPzWAYw9Qy6kd1JpbZ4l2RfYpdQ5RIA1kCskQ0hVmW0Be7YyBiQW
kw5vWOQLfRyYs/T/lTcEz67P27EiG9Ed60CYXYcIMFYvE+ie/0+Hk7Zam5LViprNRTof380fbf+7
Oi1NXxLcA5KNEI+sdRENGnSgMGzLTOp2coHlvVJDtj5MYyUixCrR1Cr2g0++iybbXlyRnLInhpjR
E6ics0htG+ie53KCCycJ8XgYwoiC/9i4SDpaqAYTylq0UuoBkgEljDTtzFGE3yY+8N+u5jGn93mD
8zuLH5EfEAQXVKUHF6PFgEKNmxiZ79PSSvGad22LaJXb7G6dAjUK6NiHwkHblo5roZcdOmE9EZOr
/h7UqzuLHn4EmytMAU7zDx+Z4sYkCBzR4B1Sq5uigyf+dofUt4Q7B01lr6wAkCrPaIeUnM5czTwL
FZktqB+h36CcVSZQNisK8bsgXyLtqKFRToBngOl2qvvwGneNm8ix5+1R2g6L3m6dSAe+nLa39Uz+
sbNTDpBEr8nsvlfyFqqy0tiDaO/udSnDKUU/ao9ziZ2cpBCmwWIvYJHnYTVqIPCWYZNPa2zS3A49
W8VJ+kvILTZO30iNX9O7HuhRlEnjdNm0N3/vdSwf89EXY1pLwQQNQaTVHYqTQ5cGefMBrG2fHxkJ
orhsqHWcPFS9RmRNi5nsCincRB+M6/yixR6/P2spIj1eb2pT9E8+tZ9rsBGtonv723aEbe2/MmT1
iFX2bN2+5ITwvPiNjSnQk3wYbtKDPjP5Uuy2xBaGSj/lSfHWrKwc7m4JFeuZC21not42MFs7PgqS
KRE7l1o7hLtFbtxDMzwL8sY+J7ljPofMmkTH6pKcOqrbWbUh0K+D48ZTLOC16eFuoxQar8o/F6zb
U17t8I9TSgW3MZHpIr1/KHt06+6RPYVGm5LYNnnMzruNKsQddaNp1ORgIuY+vcDNrROP675zjv09
nhmldOtrnopTkssmC2+NIxEeabgppybIHkULVlLzFTISOWxyOID34U1X3sOIUDuawnYYYti4BMKj
iRYyFSKTs1pssKmdElrjvMld5OFlhT2T6oN6K0DnNIdPsBJ+bQCOEpFE+oJBt6f0EVL5QSoMvNia
Y8wHxuL0Gs+6xHo42pXXPxYtEfO2BUMVLGoUEvsH1Qj3oWmg3xIPPI7yGv9gZwsNhtZ3dyoxTxru
tnP6hfk8mu50imqmIgT+sc66mAYZA5B9mmw172tskil71w/s14nGwvV0lyZlIcwCsz5Y8gQJ32XH
/ykXoNT2evPxYqikvOS9KMDworXt2Qnevd51kKUklxECJQsiFe4jY/qpO/ilho/xXquPoYwtaBUH
0TT6COfZwiHQgW39apB6EiDvJTzTyIbaLYk3nBzrlfemt/U0e13ZI1hPZUKD/sPZue2Odr62DgSP
6YBnYE2y7maCSs79LiJSdf627AVXVWoZ9ZgLWl5pDInDUmBei1n0PCKLJBY/ABcEKQJ4YK0JbuWM
lYQJFHb/01OabQdLDVbdsZgkXTQ5+InxqmP/EgZoqwLnyfWsNinlInOJMRvcCBePn4RaUOs4d+ur
rEw6wX+xQ9JwqI8pn3BHiq4PjzMIE3aLhWiiSY98dXT656sobNpPYSfoPxTOTzogGcVprWWvMZZx
SCEy8iwF0xtlhQwfK+d55sSZG84oGQCaIK/dlKNhxxN3NeeBBvoslMymzWJjaRArBvpncm7+8vrg
VHLQPMRP1E7niUe4nTU/qC8GcVD4p7bITGpTyiHixFcs8nv1pUHvDHThwTTHoWXeyDCCHPpl1Sv+
KR0Efg7V/QQMWAElKP3wL42W4amD5KZb8hhY2ghgDwPeXCbcPbo+HVJynYFFNbDPATsMgQiNZJbb
PSuwF/fmCy92OhXU+7JF/PbKNFXn/7iuIEE3NmRGL+vkkoVB18nww9/cbQS1qUemYfqzFJ0MqYgR
RZHT99OqH+Tac15KPzUwITxb8RUaITNqhnR5Ko/Cjd2TcEV5IzVaNCAOvEFccHlIxR6Y5RtpUYa6
b7UiXjUYbVJtcjZGO7k07glA4GbYAvYUJbmlLsSHIFnVWZV5jCRepZeNnzFiIzYv4PqxP00Rvoi0
Vq6CYGZj6IA/Pmaoxe3SClQVVdz2LyWW2Ik6lPOwafJsVPiSAP7Gyc9bpvO6WLAzyvqqutiGigt3
d3K2CMRzEgf+4rKjXKyUeRFij3xVhxMCMjpiSZ26DgB8KXuYUIyaq+OIG2bR9Pi5yrpkDtTKzzEf
8VhE+zYzgc6u8ohNMInR1ZwAebNSNYGJLX5wMQIUUR0g6XeCW/YoLjPZ4PS9l85hE+bGj2ihilP9
M5785N93bYvJvw/5DuR99AzKcF1Vy0nicavP1qxBhpN0qEUucEo/VSSXmIwza8EbaqboPSJxpEwK
2tIr2HIC86VoKQV0JJBSj1j38y7Gl3Vz68eUxLlXmdFECSzD7pI5bBLvXd7YQu46lGK94sRDujGk
zabVIziGnU7SQ2oHbFqkfwgod19jAMVKc+Yo6+OO6T0QUWA+3Us9xUYBc4pOxQ1Mz+ygDKuQ84Hx
67XhzGoNo0g+pscg6s5GFRPrWr4kEP60N/cVCmXa7VcPEKKJN/4ayfZ3KT7RWCEQr9hNp8QnGzPG
AgrhKJQJF8scuC5ALvNid85M5Ly5hLG2hyWnDOoaxAHlB74aojCIy1ltbdfj1cvV1dsyljTvJsKl
IKmzslLsT0uMt7B0tDGZZLn382OJrrmURckMYgo1QtI1if5ji08jBO66Qvlzo35ixl5YvhEC5Wkt
hW8urwhavkIJ8bN+y2IRqFqNZkJWcQVrOC5xm5ERdDq7rt+2GaJ+xQCUcWzj4fcO5b+R2itdr77L
P/+WWQgxMqiMNGo58bzGXd8wxb0nAnGSpQ70+ge+cb3pf5ueMseCOH9FnTdLeyP0Qu/33ILbOos9
fiSsWtGalg45dXilp0YItQxq64svO05EUZ2lPA6OXtzSXdySgDOarKIy9CeSpniOJFeia/okWxGG
W1VbBL/H6rQn3dg9lDmxBvnCj2woRqkhv5WTerb1+hYegy2H1eFbaBnmuU3Tv8C73x6Irc4m1zWG
+5TFI4IHDTU7KkXezZe2NUHaSksiaPYY609DtUPvQr1vkNmkWE/0PjX9Lx7xjTaPLIE/Ept7oB+K
l4eSkB91REJ+89E8WeGR6lSiWp7dSjK7IikGViMWr1r5GNlINjwBdYwIKwktUbr3E+fFeyIPnLlJ
rl4vpO9bRYnmhAhFIUnd6ATEt9N1sEJLDhxxquFvJvY3/t9/GxJpiiGGPXd2kzbrNIJTRRAEfbB5
fw7QkSdVuxzKmpmvWFw83Gzwpjq+ZmgeBcD455P7h5SmPSN11lvW0GVos+IHTeCuvMIKMS8hfo/M
RY4UF36KdLu4nwxBR540IePSwawC0ibnpl5b96ji
`pragma protect end_protected

// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
vFMpEn6nLRGO770dxkuZnj9GEhvM/M/bITMa5hMnLDo2XObwRZ+OzccK7gv7AH7Hd1fXjMTF0Dy0
rZoY7VX/z0GpcYJnbxvCkMMtcZqwGnAKSw/5BdDUpmiJ8nSsdobeH2zFxHFkt+e+Pd6ZyGBskyCh
gfAH7my3CvfvdCDmmGU82m5M0qm5Iz8y1CEjnAsABoks0Zr4lB9SbnxVUL4ByBiuUdfLxDrGEb3W
OPovkapI0cl8ZMfnGAUmgf4oJT5e5lfjjux8vHLfig/R2KD7dyNkJYBF0m6lvUsAGA+GDSPRvG1f
rhiVF2d/HWZsQpaSsqKIqMfsqqs/+aebneKbUQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6032)
Z9B+fLK8n9p6gr8R+qcLfqnCBfWFLtivyvTBC+cmx3EFBpf2yzj4mW13c9U/4vwEdsXA3i5rVrJ3
ymmHdLdQK8kVx+dvGWIj3XEOnI2v7MZxTlrhWj77VssAIy8+ybiIIM6/abQc47Mb61zsz5hpH127
7kU77/AKtm2H/piw66yd4Ej/Nft3fnMfqTXobCFuZ02zk95mAAhT5iHUQkLOy5J0wTioC5gVOV7q
BaWTwVrEiKhcY5XQVGksTvgkEYW0cF5CpGWneDufSmUUVcd2H7uQMWmlCY/SNAM0RwSyYlLjP+nt
NDqveDl1Oi0Ike0KeXCETnVSn1+P8TtRuUXwsi+BMtzDxApg8Rew3zCF1s7mUe3UY5l91RvPS0ex
xA7ZQyoAasfqCOgOZNXsjs77RKyD083hjSIotbJST7FhxmWU57ep6XQjHHtaM3D3TFB9Jy0D9eWj
01c96YaE4cQh5UlrJCghBQA012wjmkuW7s1ke7hW7r5Svq0XezXGXd08cRwk/XPxkB1q1xbedvPN
qw3MWB56tnfHTIR75N5qpxgOH14kL6SfvzdML4WKyjk3BtcK+YHuI1TzQN+YUYjGLg5mDfFyGJIi
pzfj21DRBma4ed/SD7JQ+Z7F1AZKl7iThtX5ZiYidvQ3mTgsT7dJyRZuIBKmG1x5NfDboA9kzboW
DqZ+B5gPIWYPmNkFSMrs+7uWgxBAoXMd128C4jBbMBZ+nmqtekkp7NLmz8SuNQ41RCgAe8cRovXC
vO3eo544CR16XXl89ONJrGwxMSdj2nh+Q1Xo/NQcAELc8JYLNDDMhpNG8yAkzAlfwYOFyZ3Mg4XT
a1h6g2Y90iAgwcfJE05QrLdt0uXyaEhBwYODRH1v6p4RJY3XMpMka6KjaX5eZhrOVKsW2FK6zkvt
J0oPbIBBKfDApq+fq2LIJVaBM/xjc9q0DBkJFH5mp39wFQ8QAEiLjIGufThyE9FouKO+B46TYb93
A1pWglTRppaGAuB0c0Hleoi2OoC9FjrRNOL+vx3iAu02+lb3RqrmWhsk4JafH86coH6t74Rclu8c
AwbXh3DLTghwV4wSNvIJ4l8U5cXG8mSowSWmRR4Bp2FWjDE5BivXVyLihMSJXIUjF70SpXYZztd9
VNt7BV6C8TradNDxpJ3NwOrS7tlMjqyt9dYoeFyGkhBWll3fNgrAojsng2anbTVBUiTAckbpp7jU
6Pdr/x87etZnvXeGLaEL12LyAdTFoyh+aMdUK0RT5zIJ5VKyvCainNYhJg519c0cUVxUYCxgA/g0
85Q8doAKkmv6MgcsDLY+uGLdOr4S6h6+SQrEwALXqK52gCY0t8qTrz3Q3bQCbeIMvLEEE4F2HqHD
asU+c1/tr2TIPjMrUOGph9WKfMWbFYM9KjxBQiwdzEG0coL4lQfUWt4BhUcbOOcWvnH7XlNFABt0
2X6IgYE1LV/fN5Fz76MCvGhQ2POEC2/lKu+9R82M2xtj//fC3FU/qssoYhRLqbuXVG9zu3JGfPlC
+XR1WFkIjcJCK93v1NR0pWZrisgorjapmffDn2GhxI30kQxX8/pqFZmS7BhkIEuAAL211PtTmSHB
nzn/5U7fnvKzoISD+r97+L+Voqj1aXgcpS7UOqYiZLJpHHgGMU/KmtregNhAFtH7ZpvNRYp7mZDx
09g7ELk3xd01l9/yHQR6Fvj1OSzolwlQXTZT66m6l1vRcV2otVH6pUp3KY2072srp53E60NxhxBX
6SZa316RLRzQOdENrWIKnE/NOyC0ArVPzKZBMyZoKG289Sne/ib0SEqfWm0sbBHr0vTccj7LirAL
deHlwSwsiU6mHv3MXNrpHyPCtsNl9Drg6wwHUqv+ja/IwYdDU/YhA8DUQ8+Od25akivBr4QzXBct
XkfVrLD32lA+h+7aou2M7Ep0sIErdoPIr1tbiG5xgV1dMOgumE+DWPcVEg5+wKILdbzAFWq8qi4F
9suxsLDP2S5j0Fn91MgoOpECsP0R+YaVl8Mt74kp1C/2SNgv9wmvPv0n/ZOrFLFbnB2NHlHyGJ/r
hCaWbSl/+CvIhL1qJ7XHYXr9JgdMlOfP76QFlOGJxM6FO4j15VscqDlY6ircNDOg6QXwzwL8CkQI
Ym312DjClWpon6ghAmvet2E1pPMPb4s3/XeQSS7khFNeQGVFOBAAWouPnnxcoMLGLA0QL5J0Dl1H
Xy97aR/BffVQkAmT/gUv25NjBRQ4YhPbVq0ZmkJKQwDYVLDl7j4jxJqkoFvgEfQcSkt80LqIg0oK
0gHoLjN7hJMxDLq7wORe5ZKMCy1HD/qcqyeqR/UXTZhpACUFO+gwNEMQELQUsy4HB/rVQIPcOQWN
N07x2q4KLzfBC+VWRN5cMj4MS+qUxtZVsfj33eQldCBeBAi5Q3wIlm6VudJ43roGsM+26Ihc10cL
7TRTiPNmJ2pworR5sAHL0wUDqBoMcjHns860FZeUX3pf9u/cVZs+lcj5YTId+g/SqUTyUGl2bj84
NR7CPygikr2P51YbLQkCJRNae2vuOm6sdaAfGFqBMJIXnEyUeVvF+LE7nW44TrNKe3FANkZcUSnX
iw9FNOfb8DV3RG1jrhks4UQKYEoNLPfL9c+KfGBXICJWiqnfv5UzeV9SoTKHctYdg1rxZ5QDqboC
ackFiNU2woNEG2RJweVJ/sYy0wUh4hwCtzf0Zwasfe/UEc8WCvhFC6xD+nlFl1NziaAe5WqeBWho
/pAL9Mm2EojAyB9f1d/Iq0plj6TwcQ1PgSeWdzy9aGVZt40x+MXK5YBM6nbRkqSY4AHga69VP4w1
GmFdO+VT+TA3z7qAE9hA+UImci6yv4WkV9UliRPU2vVnffeukfy7frQO6RgsJ2dRqOqKvkQ2uZ1W
z6EGynPHMLugVXr8z486GVdwYYdPf/BGi5DjACrnNl806PweIjOhcN4Q/xp86NSeAIAxtGA/W9n8
1gy7ongYpjUnQMSqwHhUvDBz2coWYtIsbj1WwT47vc5Ln/KXnILWiu4EDzE7PtuVg108CKRHp+Yc
N6QIXwRiuxRnE7aXpUxAWea6GggWc45fXcJ2psssRkvzdFbcvALB2CylntihFaEC6ONhrpRMvkM0
Q36tP4aOyU5ktBUVSFuRsA7E+sGF2V9yoK3y4GdwCkpEQjVIZRz7Bl+b07iEb0W6T8smjhrVcBov
tmuqQPJz9bkqG3Uon0DHINuczcZ7GrU63S+zInHcgR6ZOfBR2eB4eLPaPDNLde1/NZTYlGzaHANP
pnBmSw2Q6lPeZ9oyQmEHRjRrzxv+TNPAClNzlLGKGB+J169TTavn73VAVevOpPYtSJSKJav9o345
caypKA7XRUDKRMj19lz+6gLLv8R3nKJeNavkyrnBaeKVZ/8OfavU6wIdPIbUSxbBsIRf/eY6twQQ
UF4/V5sWmYu5rK+FTZMWAhlabEXjiKsJgTvvjPZa3nUsVOBqXvAOLyI35pmrY1Wa6mxMa4m3w6jb
I2lBQYxGp5eGazcS5r+xozYeQIvDB4Mvy4SVBt042XL0mpKPAtQdT35kECZGTnNbMh0TIEvY002n
CtomeH2oynHrCA5ZejNwuwOlrFHJDyxxayYaCraJUfzFlQX23/uopNY/GS+gXpME8t3Bh2r4jY2z
aNJdlDSN3tb2emTdI2V7mOua63jbhBYtOhsBRq3trdLKVCGN/N8Z6O2cLFjQ9aFS1Yg3JthnUA7p
b6LZunUd5fxZg/CjIoNWTz7MzZRCIpZ5b+ComM0HUVN8MMxeBdI7OsfAtmnFYj7GUx+eELFf10vt
saBHIup4mEnekiBVdQY5h6oGQfsLhOEDVHWI8BouGvlEg0ewuFz+dD5G31RWiDUReaxSi9Zdgkdx
LdTxAH82oJZkDaGn3jt25Y9z2k2cUp4D5K+zQHOgq0G5UMgWMYjr845Qpc3CGeeY3x5rPme8GVsm
J1lzgtmyCQK4z2RFSnN+kvT+B8/7l2/RkDQpq+wMnljbtNEP51MIIQB6SowUpcj6isZLqFxrc04s
JEsiNQI94+kyV/ketdvocda4YBk2IHKR0yMRDX8ZD+PV1DnUOPLWQlxQh8CyFCEbFGUWS+yUHNRy
Wid0Yhdal5cAFMb7FXORojLc/Q7TuAYTxtWuXNVKNDOLAytPkWpr309V0dL9vBlXFn5adUw0KHpJ
kUNypz7DJ7cQCQLxNNMGQhIhqKxkuW/kHHoKkX3dMFqkyjt1AyK15B45GNLYdWxFcPBuzZ34GvLZ
UE74bbSSMOQIQTnwRLT2YN7qlPmlD+9mxYs+QRQU2GL3Hnap35Z6kmGRkFD1xxhiyqdX+GagUVal
eaE+UGqcvNHlve7Mt74nBvqlz1/iXf8ta0B+/MdKrHK0RCKnHsp30ZlbuT60xjpWkECDl1WqXyfQ
mMsZvH2gIz+IzRnd1f1ALWtcew7CBnRqzFgavAiwhm98tUeme06H6QcnUTAHHVf6ofuSARYItqRq
nyuochDNGeZfzvybU4dScDQh5pjExzHoi9SpgxYsjxmrgtIN5sECqQC/Xs+m/uETQ46SST3g9kDB
YYYKxwsIMRVBEosOY3jLltYy4dij6vfxbl/Vg/R0/Hub01R/oTHn9s0nhMxIF+iqhLlVs4BB33zG
eWSOpK3EFgGtJeEjANCE+4mXcZE7TZu8WKgh6k/MaLAgkKzoCr2uaavWgnkHQFavzD0d2B4MGWiv
+IveQS4O0+93IQDWGe9TNrwI1Rx+oiigrvP1U5ms1f2p6/KO7HgfH+bft0GRriTW2hCfeg/PlN5X
aJzwYiZCZoEWCwBwUDstOLULaSgOam0mTt1LpxwmMXs6PBsIJkhIttvgqGmtAN0uf+LwhRWj7Wyk
CPjVMLfe3Mec+eDhbu8Yd0nTPn+tV3JmUbefkHufpgDw6jlChruYbrpvF2G8Fyqu0cQYIqR1s3m3
J+wmD8cXS4NKtcr/pwSxocD8Z4Cs0cFLDfYIgcg4PpBBahXVrA7hm7jAaIPytNuX7+ktJbj71hJi
2YGf539lFG1JX//rRYkGchVauEBc82Z+l7dCw44vnTeZ6i+45QZ/guuQRDuUT58+6X92YCuROewU
17doe0WeRR+MP7BjxriI6ghR98VPmIm9eCtxaPsMM5cIvUkJXTey2PB3n+ln66uz/ySTyvY4b3on
JvNFKCbIHVvn5bByU+N58FXu3KGaUH9l+maIB07JqYdrXR7TPvtnbMaKtvPNCwg1YfGd0VmZ/Uww
OM0rU+T9jTfj3+X+p+0hZKQKg/RuAJsJhFwQJdmiRpvkLjeVfMxgPQp/hH7Nk+HJu953+SWrMwgy
wD61KMaWOB7Gz6aSwkUYHQe1KQAfG/w4xw+NGOBK1IDmeicNdZquhpP3uJX6ynLyVFsWxObPXcSf
S/hzKVUT+fJMNtvlQcpZ+7BhCzgZJLC6FiTsUGvEjSDZPLvq3qwDBSniDfWBqvuELgX1QS+LoymB
lrtXH+Sy8AhS1K1OdX+rC5ETnA6J3LB1h7gg4GfJhfYtbjs7QvbTFP5NOtC2z/NC9jG9xafAcfVc
BJRYNCiXeTH22l+Zv6ZjP1ZHaQGO96XDFigSHs3XwN53X9f9NcW5JoONJtVNq7Ig8lkdGEtdAtez
me54rXSidAAlPemAQucJ1Bf8FStdfeZdvOy32+za8dyYmOeeQd/gqwMiwbUiwuuLujbzRNMDdnQ8
6KzYVvuRXZgQzCKZWlwnttrcppP1KPaPdwmrrxoAuuz9x50w6H7cdZwvGVgrxGCm/nlVq3C/Qk/E
fagaToRPH14iYX6dOdOyMe+L65HkxZxliT6OKvBYapfcplS2idlr3mqjc+3jNWScFxeiHauEN40L
cjVxwET/si9uONcW/PeCdU+fztugjr9MOUjsJnQ2vapFYr7U9wQQdVEaS6UJv8kS1jgCbpEEfqNY
05ZX5+ddYl6pl9Ux1o1beaDFAZ/wOtKO4vJiJmEGAgBLttehoKQtUdx2CZWJUzqfub1Ih4nh8SSA
UgG3JJTxOsA7yAx6QS7Po+Jn/bDi8CgRXy+pLVmWGDVk8zp6NsLvV5X9ph3nnlMyV812qjSibf05
sXa2htUKrottRTyY8MySSJ9+Xp1fV/xBtENAc3dpxv55WDpGFAnEMT+kMBkg2QgeBLDQRiqpD4Oz
ejTPqkAp0BvC5Ql5Mb+MVTA96HWJ0s4/XB7tp4kB2o6FEPFrH+sVwy89jwOWdZh5nrPgcFQVHssi
vdCWV+GhLSGQd32HfByuR0XLR1UPUaY8Sf+lJ8GLLi6JviRDuMWHGQ84jsrUNHQNvtwTJ87Rnj76
mcHx2k8PpYeuAFOI3DnTrPDxJmu5tv7/xMSihkGx7Hj4bHW8VxCxFDSjpFz4TOnnLoVYfEpjuLIo
yx0M+DHED6PZ7fDdbjM+VfgreLg6eJWaBUk1hVHqO2cZe7TciLBjLmmp9RK4hjtwqKrxqc3GcPBc
58DHrAmU4Zcnb8lKh7FVVyVuLJxrXUNXN9HS2ThSBFIsFXmH6yVOC8vAwhQgP5ejIXaBLI825pY3
c0UXX6f/DI757BGoJ4skJQU78i7426VHQbzQdiRa0JZZlaflnnzsWtVxTYFx3E9Rx91i5bi2Y98R
318WFtZt7qLMbD8AHGki9CeMMWeBzEBLuQ/exikcZw2zGW+2FWQU6ovbKHirhaz/n6LUFO53uRjz
uzItSzXDM38CAyVzn/MDgXDzf1d0pdyuIyyGqfNOaOnwmOeqXVTTfkV1ZASOQuVheilvX7OpE2yZ
5Y1wsdqs3qOrWm0uV/zTz87WuebzaIJnswj5fxhRNv2QKeNyITSgirR2+yUQ/vsQVW5UeL90HDqq
C3QnCprHXkYrCe8riqy4p0h81SVJZF7cMEsWb2pa6Qte4yLKMx9oIm2i18+sb6+4p/ocf+mOKUaf
v3VAufkk94OYX5O/mxhKlB4pa7ieH28dH2Old5YcSeId4dGoe2oQotn6wFaxm+/lYdK6B9pHIOz+
V4Ro7XsuF+5Itsfk1R4QDoDGthlwkKYrWJyczOvD9gxyj96sVYWSwXpNO5+HLHD3y4TrcNtBlLsv
h2d+Lxw5Rv7k+LD4D7nvjXkPHgMsYr02KdU9bcfkSDkd/y1PTY4whI3ROuwozz5iyXeo1eSelie7
cXNKa5jlLo0LTNq/gg/m0SVUPvVqkIKBXi2SA4fXAQnA5WR0Pn+AFGGo3T7aAqOGl9+EqqQupO50
7iBm09XR4Z2bLdRDom5seIVnJvub1nOjlMekXXZqYCx3p33Vx56QMLvDBzcOLhVczMT/vl3ZIS4J
jNTc1ulgfNIZT9t+1tPp2giJwKtdBmJyzb9z1zto/q+6UTJOAw2nG0TbiObOotHvOPhx2iVsupDI
Hg8ZqS3uN/ed0LuGsGmI99RLc3ondIhmQcjtZ+ihvkYvD2uLe6hj+vgFVpp4+Ytay2WrLc2SimPX
zAcDD4LrW+++x2AxriD76Q6FYFjzSed9yLt/p/3uhLvJlrQNN+nhCPsFKYZ8rPp4Z9a06uMazRoM
OdiTwWyxPSSWx5kqeS5zAY/c1vP8bVu4J2FczD4Oi7gcqnbTxeNZV1f6Ju1Off0eoZIrHjDbYjxf
k56DkdJw1lKYZvtTE1JnRVhFrNSFUsdktyPA9+IbrHGKPoLkNUBTrt8HMSwJEK4cPNPjcK97hrOr
gE2z8TS+yjuTgVWcyzquNn7lgUPQv1l0iNolUGZnJc0F/Ua5BPM83lyF19CtEKlxilm+v97Lg/d8
Wn3hRy8Wqhjzan0V++LihzFDDu2OYx1aGzlWpiOylQiKINt3OQK8AI1fOKeqp4uCMqQpBDw2Y44t
DLLAMS+Fv7+WKasCdpCfp3WCbXWDymBh2LDNa7X3RNAnOklerTNQvBUIlLdg7y5zoTrto8AE8+Ug
CZwjlRXnS88wUvdhr+GRkIxgF68YRDEUZrnPMCgFXXVjZe6h0vwD0xD0MihkwW4aGR2jwF7/WePw
jZmCjuSQihMMEVfzkVEZm+7qk8ehup4A8TMDYd0ps5M3rFBHZeo6/1uFOFxYJfI=
`pragma protect end_protected

// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
XHHrc+D0970YSXsQyWN61cxCWgkiIlOPtWraaNqJTg/hUWHlUtA6nLH6C//YQ3UJWgUWbOZIEZai
GRtJCKklmRkGqIclLBpPdSwb54gHSvPS9i+RlmWc1Ft2BGSsgPMG+Edc/F3pE070V10HK3RsC9nk
sK20QpVxPKPM+ZYUVriVmy5xVphAPr0YD0B+1CJTzzR5SIz/vthqZGErYoBIJ6HY4+tLQf9BoCQy
5pXVLXdhpx2NLvi8pdD6Cun9zgQg9d8in51I61XwikkOEOc9SWTFUY9Yn0T90ltGj+YiX1NNMm3e
fHcUQYweft5YzcX1M1Uv/DqZDZ7pxBceaK66lQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 31680)
C4VyRIbV3pvEGwmN/mEqJLIDiLyfD8sQYx3GlTEWcCgLWNCDIjMki2xiTx/5DAYjjcoZMeRLaQeJ
MlOfd5WPiNoed2MmjhDFdLDZdufR46fkR2f3znrH6HPuyo83zFsMfIa0ajCCctLVIePZsl3o6rq6
Tf5A5wgPvDCEhC1hHOAAao5sDKfNjhwjDiC3Jt1evpYoWyc02dtBPpDjqukRJ5s/1f2S8IXEe8vm
yxPZ7WYlehDwBgaJMD48gwyHmKp1OCWfhPFg3YcZNlL2t21MciE9q6G5tKD0YdryXWjOTVRm+Lsm
CPBHN56Ab3Dja6WX7k8ZyZEA5cjcJCQAdJ6bxOfUhO6sedg079AJ57H26EkfhAGQjeOCjkFKDABi
9rdLczKO/Wi10KxP/A9O2GR73EhlWeJHh2ZQPjvtT/V074s8+9iCRhZL66JKpMp6OXQ3pApMpi+1
A5WidURbkDIfNgl7607S9w7R4GisJd8b/GNHjdcn9/Q4N8yZy2fMScgRkt9uk4ouLJpw3z/vjvvT
q8lU+nDJ+H2/Hst4iaw1csFgju1biNPmr5KnU7CV+r97nu7u/UymRDNKxfA1TnUbb7PTtchLUBHt
8wC6p2sdSO5CTelaHfqBdDrfTR7L3/eU84tIoazfbUw94EfO+RSA/7CL5AwA2P4lkEp8LgJVez3o
8PY5Fo9dV4rkJzuQdB+boHf8y23cngfWoERXyUmQzpbGv3RwKccU4xinhJTbEFRRRtsptAwhH1eE
GYkKuTjYaAKaX8Tr7b0qq3jVC0BsvOnMZZciXAv12S/l4Wl7VKHMAlWTyYXjV6un4fF8i0rZNVSm
UmSDefiEa/suiFmHTjgVimDRVkyH0uLL97XM3gp8UzS1dvmQrbUAEVkgrafBdwaFkUhnTeH6KCUZ
f929wYs5IFuvIVdGMa0Of5K8sqHWQYdr93fyQwdccRyC9T8Gn4+SUC+vK0eMQJvOP8X5L0iOzj4L
hsAodlp2/sQIvZq6Hy98iGEBagmaIIJVJbiUWSk04gAuV3okcaHkdxJPeeM2aR7674+6MXsVU1Yt
dMbUafA5KSvxeNm51pd/vexkq6mR40Dx+lG5vvmIGDGpFMVwERGbFQ+yym15X/gywOGcgd2Vt/jV
b+HBxfP8+f2/w34M7W5uFtJ+9i2HvGpaIjEishbP5zi8GXu3EmdVPC/U2I5tWnkvLUvEgQ8/jvV9
K/khDCIOB6Q3LG7GOfpKVXKGv6lb2A56+Iqysx1Oy5DrLNve0swbn28ahkFZHmbkKn66VWz+LdWt
tHlqe1nwObjIrT81UJ3bvQkOoXKWLcwEydekePajulnZHHJOKEs//Tc1Jif7fbVo0IpxzYWzrbpl
r1tIENj7AgoLi/LJ/r5ERlAKvCDSC+sTsA1FdqRY+LFUrgDRybri4ssOvgB9E3zjZXhTO3q98fNa
3XD/RMlGp6U64TLji7ZCbwmr43jEBYx+15f/iiFd1+RGeIM42ZiIXZLTJGXA9eN3kuIE6JX677LA
sQW+XLh7nK0LSypT+iiKRiRProLrnIk4AVjSN3SmclNqVenhzxC6yp2hC3blRoNll9uc/w9CCGV3
11AapWktG64oEEKhcXOHmvN6GW0CKpchePfVXpOiwYqRJm4DNXQR/5qPTAagwC8lR5dZnOCpUGpY
pihIaRuGbjbg/ZBk7Mb9wXjUYLqJ23KO9YlVkTekhqERzTX8ra3t5LOAucNUixyx0Vfeaf1gSkhm
xDUD0qnZdN4VAsUccgarXXz0CGzf11fBZgBOdQCZPQjb0XLNwf4LsiWlosX/VusJ52NPvREZQAbr
4KZa24a1SNImXvMNprTo3FpNyNsb1ZAzArtQxujd/Vc63isBtH+RhY6mN4SgEL+5L6jr+WxTyleW
LaiN7ElEpSrgFVQ3RUYhGdb9PpwSDas45iQM8k3EBUJEwLqpwzQnZeedd1GvxKG8G9QXAhK6G0Hv
xIa9v1lJ0wi5WuV0TesD/ye/EAVzOsLAhulCoGZveDeFBmCkqb3dAqFxszgP85x+1nzMuDex76l2
rpnuPokJwNsE89JhrA+rUOjo+P0TLWWM46cN5XvtRUd2aKfs4tecLu5/2EpuA9ag3x7MsHcgN01W
u1CKuuGuTgj1mIx0dvqqzYsDx6Yev1jkqBn7fNaMtXiRbKDgtev1XoZV85nrhtn9I9pi//7wDaPs
2G0AhRD7u3ZFEGYIKPf2vGVK8q5Q53nH/sE/ySGFvvwt9YCaT0PYqi3g4erI/es802WM8x9E3GyI
HPCb4wZrWHmhflb5qnWnIphdBMJJde5N4SL6qpItc9/ivXyx/ZTsrd9mLOHboG+LxGAg59cgTna3
y5joFW1wQ6ZEZWzkDNs0M1TTUbG9PmOR9hYEzVdjSzE6zJTxNxY8CBRPeaMdQbLyDA5vjxEtzDT9
gdJrkvhFGOhsR//SHHd83cU0EkogwFgkLwRrCxT/FZ22dKTHxGYE2UJNpQN0HS2VEWe4NBguJqZZ
Mg+GAOp5Ouf/TWSqhD3pvrvfy90mcDP1ut+RGgUe+v1NElYYDayYO0p5vjz0pdzCV4avZn1N6kup
K9THHEwPQPCcxsnZbOVIU/hbAZq79sl+CxeHsLNc4/8ytFOHjgn3t6aeXSA2qIDHy6rIZL1uZ64u
msKuaVjCO83+wxZfrMvguZwc23jyAMYMNX3E5Ckz8GmQncQaRdexOlOBVCnbGfyOm1oIUxKZwwIU
A6PmpoQDQyGUOwjFMbSUMIl/vOoRplk4/7NRUSU5aDlfzGOXOkts/YQDJ01xtVwysRkrPdJRDa44
83OY8PLBxH7C0hakmTYwv+k4QwlTDDDFUdpBaZhlfsfLI0yi0ER5TWtrsdkkwzIVmTAxhAT2TjOs
WrUOuLoX4GkBG1bsm6ifoL3OuIcNK5i6syUaiSaZw7dtu/l0FwXrJYeSYn7qxbU2xGyhtTegkZwG
j8nPP7xGcBk9cCkL94/mv4/hgA3pdgyApHT0S9Ere1zQiAjV0cfII2Sblxzxd7bX8qK9Hf7I/SCt
n6wdOLMU1e+t0zIPo6WbrYNzPsdyWPzkg5qNMPy7lAOh1Gv5CV2GjN02WP0Np5fV1ovodFbvvMjE
/9ohtzlR8BlO29hs98zA5B9PCB+Uv9HeGc9/BcEzrdD//1C5hACbhq6hEsaX1DUi2PSPqdgNJyYX
GH7cKBH1c4zF0pM+t9lQeNNFlGp+UjcQKdeAolfX49LZHGEYm9pt/gGlxf7crSB8Bp2D2eHeMORI
AIx8g5EDMRidXeDPlfZXcsTU4P39iwrz9+whEfZBIRNa/xOqqJBBUm5IkwIeQFD4BwhH5IAFOF8p
BHqudO9JrZBcQzFmZ5pA08JuHMNicqoZbfzS6UFJGK8+pA07CoFRqGQ/cb0+qUK81tBk0jeLwXbG
9ln56QMBcUrtMICk3Uaom5tplvmva6iH28VUPz88dzp2gmNRKrq/IiSMo8FUJH4/WjHj2nCDijan
Vf+hEM0eWtMN1YyQ1ZVE2wV2fKum7hixzSiXVPBBLTAQNRUVlTRxp2yrj/dPKCI6/SywzJdWlJVs
2S2reJmcntzhXIbe8tz9LE61FKnOEWVB9ASwi8MVIB0/MfQZyAdPt+OOgAwJ0MJMBb7DXzylebYV
P/Q+fQ1GzjLeo0yMUJftiMgYlLXM5LMupowTxHVVBh/3vlj15mCCc7sqM+hCf14FaDbqD7nSbbXP
LNQerJ0SICcl5hgdsYrA9JNUXyNLs+USqiccQ77Lcp6+GhLqguUDAEnXXX2z48ZzpxufEFjrf454
UAQyq3v3/4FtOypEOmrJhGkhmST3m1jnSENThm+R59Lna87wqASjxQKwnyeh+HWYWjNbDyzOK6FA
p4S/D9W8BSs3moEW2YEmLpfYaU+S3b8ZErVL0CtRGZB7+wjJU4jbHhzajYoRWBZbUkQttVV72A1C
ZK0D0c08EFdRfHc6Q8KyrofGBQxbMFGqYFBspm99lv5aL4tbJLLuap1CALcpWnEvc5vcLyENooFg
TTqWvo51SnmZJgXx6ZGBYt9dXCKzOmvXgBwzFjjPlTUZ6NhIAPfHHJUxphkkk34thsIba0bUF2YY
AcvshdnC5BPwIrGrDh8P6/UqYOMNip+KPC7/Sn1gq9dnx6XpUM6lnNFjTr5DpL7qnNUmNPK9vbuG
SgfQzVLg+3B3t+ZkwGGLvd7yBJYjhBKnD+WUxSYVTalT7zu69TuLp53yChc9+f7guH0PRkJlvHkT
oQbT6SlOn5/ceKcXls4r2iJBr3rinQheM2cUMt6faWnEb5BL1V5zzfjxpapaZzEoUl3RA0f5xAEe
jqHWMa9sQkN9GV4jPTIzom2cluPPdVOfgRh6H2CYF7HYlA9Ps62/0HYjsC1CQziGLRFyHdaqBloG
tZ0mjbaeFJ51QxdVRpfYuJv90LBgPGoC730GzqMQXKTDgjQMleOD36fTA3JbAZXTZ0Vp8L151h3t
wztYx6UUYvtddh2jTwqq/Qdb/ewqLWADB6ZrknO8CO5tNyni38EJjXmbUnA3m/E680ZvXGtTPPBZ
Az2lghuu7Azyn5/TqoDH31nLqx3MJQPhfv7qqoqWoP4tcWQvfyrBUzEZ7KUNxeHp/Q5+hLNOwjpf
H7cnSRPzgKTHhvCKWdheH/BHs7sShxStRFWb9c7iahKYRItesfSA0ea0+g8yy5xVdlxwWwPdxU1q
hSpEBqr1OXjM1Fm7NTb5ktRgJ1PplkSw4cFmUf0540iKeaqgAy+xIbHqmEumm9cQ3W7cbXY7egpD
gtaqNdbSqWoBmtHldblT+5Aham3Ru33Ty8Flua7h2VTZ/+DntpzveAANdmNeye504y3R+0bjvtS7
Hp/+SJNG89FuCKUMM0kia2TL3zER5eaF/h+F5DTJTDQsNWhb3kxRDfclh2KSaxv7Rh7jhHK+/vJg
nl/9KQDRTFbFv2fWw8cPHabS7587UrR5Kp1d+u/9i0E0C9V0zFobLZ3obRSw91J8zSZ+JOV/NGrr
OGVetl0ucwxReHrPoErJdlauFpO+9MZGT1R6wC1aMcKOP9eU5jSxGQbVpH4ikoLjvl72mcLw083J
GKKKZuQtz77UAEPfe1OI2jpPZyiMcaZdoWY158T1baGRWOEd3MPvzPZc3EoHJxNJgr5KmfUpN3Pl
6uoRl2ZdMtNWwb1k8BG3q/7wyeU4Z1gcct9hWqvHqPA3gv7YVivQWmlqMxqbq6tg1uMNSuKaPdQ6
stRu1h7ZLam/1Ebhj7l8+qsQ1I29h+KG2gNMVmoberJmfcvuS1e3C2h2IZ/qoOrwwPvUSL3p+JS6
+OXyG81zdGzB/wzNA4iUv1sn8j33aBoaPgPX9lyw9kr+CWhrqONdSKTU1j/tj5g+vcczy/L9Io82
i0KV77h9OXBrg/xYgOfBkdYBuAa5OwgRo1L8L6m/T2Bc4SEn1JQ7a7Q8/LEAQVfIS6aEL+eUK5jE
zOOIE8BFxw5JJEExNPLHZVWK923pFAHSRxscXCOfAHKXLs1Jo3n+yxAgVYvqg6NJulCEkOqeb4T1
QOaamOUT+DaSXbGGF/fLzRIn1KXry4oKyi7b4PICYXWB+NKfmsc5H+Hm3GH8ms2C34tbYrBHq6nW
B/BSZqGnL7FwqKWvllZic5ZH/B6VHDICew4Bn+67LQWkbS+bjqZK95jyGuY5gpRs04OAYaH/ov1K
Z+b3uEAMtyF1P5qWru2Q8CbDkpI8zprh5fv4zlB/AqFeIhOq0fezf2TMCUd87R84XwsqJVlb4ltu
yenxJMlYUPrAY82CfUrrW02MFTNqeLZ2IXo32mSjk6Mh7fCyqGXaVCakqR7Tbh0r6F+MtCXloHu5
geqV/SabCv08z//Pqv5MyiPuk9PQnsuI4l6+0E7EFUwMgrftMKvUJMnP/jP4JRZHAfGU4V/pMfAZ
kNCokn8w9CRmJmU63mSawDT/wxjqaV6e3vYIkK0rseUedzTsBadduiJ4MhUn6FtBUVxB8qExf+MZ
Zn7DpPs48o1vBjYhtZ+csjxYrKPZUMjHpX6GjjT7LqMbBlWQtqPILtJmEHo+YWxOMtctYUbcggXy
Pgtgf4Js3Tr8/zgLIVCOa98HQULunl/VOxoQHtSRiP9pq4l2TL0xFIAnT18SPiGC0Lw4YatVRyFe
KpG1RvF9r4+7cx0I1g/DgJzi4RI1ysiNM7xSblKfIGOl9zjy/xK/cdIo9+EhKb0loX6iYP4eOOOz
BsYOCwYsq9lMZ+TXBTcbyLJfVYaEAnrwxR+kMhE+qX4pa9EhZk2GTgNgnDTnkW5KP2udDakczaZF
bV6JDyEDutYMcF6fHGs/LkAp0VAbH9RngM9yLUAP0kilmQhc0yKIZiEfSZU6XB3BmukfgT3VRSTe
Gk5bexpWfvtm3tyg0+TXGlSuefZDy940pDWLb1WeZeknukolsK1bW+P4cC7hQvwXhZjk8x0t3L2B
iO0m/3GIYatYeY9pXD76exA0Hn+wFX8kKiUU4MtpbepG2WF7TtuuXNQW/KOL/Drru8i7/17S2z4d
X2so5EPd0/SJfit/jlidNMvy9eGI7kzIcf+iE8NG9PywqqkTIcdzIUtqk0l7arL82gDWkQeWbSLc
3ePJ4yVovjfykizhWgBeeeEQ/Y6dFPzOWoaqPNvWHv6MZqvhP0laTYXlWMsjEZj6FUFfp9CQYPaA
QoH51Gv689e3VB7TOMxfyrhixVGMnxQaVPhDENMV435M5/lgFAmqNyKx2neJHZgRD/BpvIuW93d8
vEXwks8HNclbgIBlG9rZdwgFwnWnQrZHLGOLrpkKiCM94OaGqR8O85vvLroRGacZSPFM95uFA7VK
8OpHvHl4+PGIxy9ujblTEm9jSBHn3PnWEhJ10Z/pno1e/HRMJJvxdFdgZBj7qFN2N2zfGQB8VxEq
oexdENEpFAI4hsGsB5Ok+fVucJtnPkHb4fVy4kLeEMLXLOPvuK4jV91Q3hagV61xlwdYhrfFyEEj
ftlNxwK0BvgQbieSK7vrEWdN35aNXLyZd6MB0+vk69H7vy8GRLJmyjgPT85nake5Avnf4eYnMC/h
3dbgdmpSlZ17GYXjKB19PuvuP/oaxbhgF6EsylTR6dBr/kgHtXShjIlXxkAUk+5XNDbXRzB+EqU2
MHDBE5vFehTQjpTGAaXLa/twfrKs9/rQstjgGoBV6u48Pt16clkZ5jbxfes2rlvTpp62On14So/1
cMHlWof6sv0fuje2DS53JqyHZt1EjlNjMFyHgeZ9NVnwUzRNKfm0Gis9ng1IusZMUxgMg/DjXM6o
HS64rV6MZEZn0HPD9MJAMwi+x90wSb0LGxLGOPvWbr8Aca/iRf0o1mkCpFc7qJLz1TytxDnwMPo9
r5Lvy36N93hYsOJb/VhdmljQJc9vzw1nB4YxQEKzCx5xW0u33lgDO2NnpTqGMSkyF4moLLoUDB5G
rDuZVRR/gck7g6XyiWGAS7oABiIlQkvOjdlxr539uNAjWtEzkenYNSITWyrcppaF5QoDlhduRQEq
Zi3UYkCfybqxmQq5JWIIqdPBIHhTJ7V8dlTfTm861syOHbwFN6v25gkZXARmgy6d3wBXvoqTTY/f
3Kng3TAtNOfTJdCVzGeGLPqyabLupH9yLeF/x5qxEnNTko4d5o+Ue8h6QPLWj7jSQR1rKw4u/r3z
D0bZdLOIX92M3tzaQSdLl+XvR62Yd/cE1YRRFdFYus1SIbHecHtOnyf3U5M4pF8OcFGkgNH4wccR
LlZDvK9SKDNpQDSiQ88FHT9fbCpx0guTxO1vqEiulBJOxg0CoRDAXmOYoqmOsBEqmQMsQzQfv19r
fXRLt2rFaTl/x9DsivxTC3WDLXF5J+yyh4HKfyTTlGAxFmQdj09jALkqFJ/GbBMBuXSyZi1t3RKf
ggD3Cf2RG0NLtLdwTWPICaAj76TtWOuQfGzDub7j+j0ni31hzZ0Ek0sMqC8gM/1zNDqMPrCyvybO
ybOnWBVYA7eyWO7ZUVOxudBwAnNalvPhuwbD2NCEVTtb/6jkEYNiOclpHsWuV9Cce1+CDd88EHZf
divWI4Bkumc25ovZndGPCS/vfhxCNt8DqncX7+MCNOod/mFrQ99kcQMe5Wf3AS7j4FJItr7fgRU4
O7UTBml9NQzUJ4TBRO5V1ejuP3lkMk1U8tIqtM0Gji8S7w49yJbXp66B6J9zurspHZyRLmKd7I/H
gt1t/DHUvWhW0cwQMuP1U5wTAhMSq1ijSH6Un3JiV25LW8AwOV0Vbnozl4ZnGqM8v3PK+Pq9R2rR
AOdlppmjIUIq6mbdn0+5MD2zHrKM1U7lDeeRXzfOp5ZWDaLIHyi3HLVk/mRqA8BzYtFF1NXDmA5n
CRNeR9rX/6FV+O/10V2P1qDGSXLdTnZPkcJ9tdgwADlwBC/ZVDO0yhPHZ9ZxjulIYSKFEfk8KS9t
dUpwAZGMFdHELBBMvqywY8y8aP0pFCfFdRZqvx6yndXyXIfjiJWiLYJDBLg3Qn+LY9A4npTcnLyL
ZiGD/P85X8vi8T4LiZXZkiifPdEA3rBi0gkgG+S+L0QaLabjCVS7z7i+T3dNfRsLjaZai7SU5RsR
Gxvm0XRw+jCaT+zr6fTOcYtJp50NvttaKEgghWC3VRAruY0SbtI2xcB5temPdKKSUEdVYhqLoEew
YD4CI/uTfqq7eCuvs6Hqg0KgA/zQpV26NpO/zZcbnYipYCAZTiqJRr+4GM/4BmYoGbT50JIvKx52
ia7uMY1cJvh5sUYWHkFNS987b4sg0IIcyBhjQm7mNHE1TiLrR+k3T5LJxwlmRO3Znc669SesGaD3
2QdouRlDYMAdMxt3UKwr0WT2k5hxjUy34BYXWsffam32KQ1esToSWSUDtL5KE9RA2h394bovaZ2+
oGeMcxK6kb+oOi3bnoTPifhoU+7fOA5ivVluaPdIESnSPkxeMOc4mGqzKdx8mcGJsIih4jWsEJRE
CLsXEXULxEI9P1/f08KHfXq45+y9eDb4OiYgC6WFjgXScqkU9vaMQTMP8quePLrw29VJ9ffOKWeX
JxgYJRrdXU2YMKmwko3ukqUrskG9S8BUAJ9MpCYXGSG5Lr8eiAYJC9keBYI5D/hGhQluDkYFolfV
Tlo7wiMHP7eN4oKwPczqdEdU+TBjqjJ7k1m6RguRw+tSgLHB6bH/Yidr2Ji9eQ74bAjd6tjA9PaC
Ez5I5qgEelgF0URmwtBTfWmTQ4z/CW4a3ENoxNECf4OeOy8qxGbZnq7dNA+9eooTNQ/7/fXIY5xQ
+pJ+jJjRbJS/QvNlJmSVOOHFpTWbgsWCFguwqDk9QrgNgrShcr/1UiQaKx9oMsjtrMEjypz14LqP
8AFKgM1Ky7nhIlxwTiNMGuFOVcMV5+hh9eRxQxGB5d45FUxthca4mX97hevvUeu2Bi5yqjNvR93w
yOArmFMfJQxtH+x/dyY3uFVS2GJEH3JqIX0rGFjQN4Y1V4Vp7uJxuIBkktYcUj3YojI43QEGD+12
EtqF+pc2V2TsPM8QUi4vxu3/dyTj+nZ6OkxUReC5zAwIszdOOujGcGZs2UHTD9vW85ws/W5Yfgx2
n99pNykm0uFYaElvJXrpKxk5sBTWntaBe1DKIvmptIGfMZtGGeoS/4jhWjYJEOaCN2hr1BEAo/sW
yGunBEwUJpwyd2Ph2bZ3j7/scPZlwtMsV3zUsWwe/nGTPNRcesDtudqH+85I7vgONnfe/vg2rn12
3Q5os7YQsmwkdO9WMK32RuJ2VlMwAZdRvGSnhhTwTblnaXhS3TqQBd9ZtYM0faqAqku5dB0klrJ6
1V0zMknViGPDTHBr19IiKeK9eaL3IyOqH4AS7A2cKIHCkonXxFgfhRwa3GXc+wKIwt+HoHgeo6AP
NBAovVLke+2ZoI/7g4677njpoHbo6gQN/JJstkn8CRzNRBO5l43nM6JF2zEJboH0tkoNULG92RUw
7zdBO6bGUofKv65Asv1gGcQasGtuEkrcPBPcsg0/OpwyVqdy/aFieAxBTtewXlRvTr17Qv/G7ppP
JZiO1a2pwlHu/KDdn+MYA9YevvOebdKLHQ/xcJCTYPR248atDS7sYvrp+jujLXnnANA8vzrKmmlx
INHYZizYtlJfBXSyp1mZ/PvfkJRT1m5DKdNAZa35W3BR5cTpKR+wHWGobTDkLLXmi6oD2jGWhDl+
nsrAiHzQlzik/EOOz/N1VJUocjkxFGImTmMSfwWKcnha60qItIPnh8YA7TpqdTHqbOaFbkeNtgeU
g+UV+0XVYntFo97NYP+kh7oeOIvNcyxLWCFi+1oRdpXXMNtSJ2e77oClr9TqcXTYc9TfoAWrYpWi
EFQb6UIW2fF0zGYPmsO2RP8EFmRVRG5r7nHCqpavr5Brw2AocecBArAKR6m8fNBQApWRr4uldhlx
n46wOK1BSZ02HLVI/wKUAQXOy1uO29YyS4bgClwlmv4BkUhoDdXiSDJc9mtjxHwQKJvENHmVdYMO
I4LTdpCx+bhtkpOwXUOwxAGH4xKJDFH0TVf00EFai5RpmtPWm2+Wprhx3S3OUCs96jKRztEXXDZq
jiEsa60PrtbPbEvDpk6QHV2ueqZwsDfAYfYUxiEHW1eUbtA7DYbZmb/CtyIqe2aWVc9TgqkZg4mY
pWzxigN+NjfuGBpU/Mtf+o//LwZfoNQ6fxr2Yh8f4IB6a5kItIqgj4q1H4Vd7MvNnbFJQyziD7cW
Rzkt5vyZ1ryDkjS0SJRWxkfCtJvfHpze44xpVT4Uz/ioCJIYMSkMQhBHsEsqc62RMip0Kl2N9PzD
9E3RpeN0E2pXZvAjfvcgmSkMRsxqNh29wTe+4QLLYBFzuJ0I2bTCsfdJYY76r+J20ELScqYCfs7j
reKorPGYYZetLBR0JZtjxgLlUFc/tVcEuDCS10mBAnxV1pKR5+vrcPe1Pmam4Z8KtLggql6mymRV
XnKU3li34gyz97uuzklL3uVRWXAljX7N+1ECIO1Hap1nNHwfYxtiCTcQDZQGcuowiI4Xvo3LEwbK
bZgqVWYg6ywNv65RPG26LQDuITnW4x1UvKi88xUj8Bbz//oXsGCrxobg69EDWkhpeQ5wMRUqg/nh
Qml7F0rMs0aNouwhlk+x0w9nJibrSSAEuzbQv68PDgJjugk6WLdswbE8OveZj954+6pUGcpaSolk
XonA1lzeZdD2WJN2soCb1Q14DFEdLe4FYAm4PkLA2lj+xIILRwFCy8/I/l9GtBugTsbp2+KhGCna
KDGchvJT0B2+bWJnX/VS4mQ3KKSc4nz+3gw/EuIAEcYgPX9IqNN2BnlWRLqrN+MbqqnoUaMMIavP
PX2r/AcTWo6ysf+KCLkOwykLyThvtY4VbRIVxqOqAM1YyZ6sGof++aRDCiDLxE3Knnq2AOKzsFKL
o/chqsm+RCRdGmi/HzN9a7WwbvFis+SNcNNPEPB30FQ0OM16SEV66ENgPggClYjKr7rSPArKIFCc
JKkigJgb7FSMZqrOayaWO7RT+byNK2FBQMWotmuWKHp1HYqIf9ygtPGeEGHBKugBlXAllpvoP8Vq
DavTYEprcoMjlCc1JSOVefGkNgwzzJAmIrYd/z/UXik9Ly3EO0fAcW4+LQJrKVzIVCgXko/+7xpd
l1Cr5+aucNGoJpXSrv7ZMGn4wG7bQ32iNq7qyY20hZBtJue1WJ5myOcFi/GJ0ZUP9eI6+rjcwzoC
FMy5fqvJcOjF2xlnstAocyHn6Iw+5Sbc0sm3Q5mHI9J2Ac5hsdhnIzJYQgwEdW3AMrx51TnguRKw
/ZiyI/tzuwDBkQWE9PbS5k61xhzy3SEQ6H6y4TGSEUiYY+pZvrbTdDO5XEWjMWbOXa7zkbAK39Lq
OJfnCYH75aBCIAQgSTLjOKzV8ih3kv2dFfmnRWAYUYdlHW0lTSTwCYCce5c+x6yfAuYVyijfiHkN
3/yR15cIF0yBkG3606uTvFP8NEOsRJbzwHwjlPqks1v3Dl5PZdwJAKuHunfRoqVWSrbhm4FaSwJc
Cuz8e/RWMlOJvvjmF8xZbau8j8k0W1gqY6NdbG+DIPBNa7j6x//ZXXHZOxyW3VAoghJTogvlZWn8
WUkGFapV/hwZGMb3YE2+0MrMNqlL4d5Sl1OD1+euVgcGBT6CzD5e9rKLcwvd8lLP8KsqCb5DHI2T
RPQ0AY+gOwjevlr2z0myt5Pa8l9uKFX80OwRXf/2o8PoeiZw4GSiZMU9YZLBT/wmEjmVExFvTzkQ
DBvrv903aN/ka6pEl2tRH252q/X+XH4hiTzB7v4s/vLGjqphQl7bfpu/z7OJ1lz4QANiw+LMIc4M
arPvXI1rsmdizpN7I6306yy3s2P1My4sSmdSU7FhBM+yIKCIf68VosKsz8cEpR5rHePPZ4VVHUcd
LsV+Do/A9C1lNahgRIAqKZG28p9XF5B+IqRseNWSzZsJfQfv42SFphqw/avfX2Hmw3/BpgGch8zp
tt0UaiyTrKAo5rvRZj7YlUT3vYsrs6MqzWHvsBJ4YsXVttQ/rv0L2OcXk07fl+pZnYqjhbEn5NKC
dgHgsW2n5wklYjb/sdYVyFn0SL7/E7OsdN4VXuHXTlMHfLgzZdCd5u0ybbDMBKPA7BdVAbEO8bI0
p0UKFViRvllPeCp4nPEbwqNGCZ3CfO/AIYo6X1aHj8fuHi8jvbHwxy+1nWg3SC9ayXNGFEc1p/vT
e9WqI7B5XournPXCI3kEy3kMjyDTc9w/7FzFccYhmKdZkLp0F16aWQpjJ7kx285BjJPLGB7tfymj
uLRljXX3hfeYqOE3RY7MJ7eB373y6LEV2jLkJh+fWAYDieDHv1fx2kCyulydsAuc8JgFFyA8QSV7
vlJSmBYMKPjqypx/CioJGq2YpB4qKK9IxZR8765IDty9RaZpM7vX2OlwGivOzRZHcQhkkhA7RG8S
bI4cJnHf+cSJL5a0KF8Omx6RG8r9K+v34dZ3jf/ja69HpqHMDF/Fcdekwged+BXQRN1pel5sb7uH
stppCf2DdC8UFWB4zLUGKy7kxkUJOibjXAzhQeOZoqMGTp0i77biVr4AflN3kIYUGWhqsg+01jta
O1JbY2U17cJgydCeoMGO/8vACzhvPDV7SbdSUW0en97PXdh724bX7THn70EC0o+xf9aeEAb+a9x2
gdsUEDVHzfj5yh0y565hjrVVrkHYUp0C3RwvXiyRORT+N1PSQszXaimW9B3qxMpWdLQOVFLjaskb
Q+x+zNyJ0knJRbLObw0tXpQfuJ3MwTG1U8z/D++pRkCTmRBGTsc0b/ET4A0vEu0fOJMAEcW9Hniy
ced6F2UDZ818GGwAMZbA9RT8tYmj8ygV2pX4l282hyxAhM3xzlnamh0tRnn7cdr1PtfsncaSmZdn
yIjYZpPLhzVVUX0Keiru/EFkjU55GooOxCKtnrqUwl1lboqFqfTDW/KLo4PDYa7YfdHvPAAyR2+S
zvMhaf/pIpLr8x8eqJH2LfPOmBv4VWbKWmXTovEXD4hlADBFO9OVqGHO0JflgzaI3CYfcYzIfOfg
qXiYR4e91FzQLODQekA/zZBW64VsdfGoRP8fc36w2EhzatMI5G0kHAsMurC043AWcHk3HQq8NE5p
f6ziSiFARDl3UFUOjT63Dg9eT8KL3lWMesxxWLD80QXjTw7OOB0PDmAdmG1X1WoLv6ZHcQk5wfs7
ZNOomxMuc8m9RwfBUvSFgcXO4Qqag/w3NzSHFIgunCXgpGcdG3Zo1UnxIlIWwzHoSdQJDv8U6qbf
TGj0z16HPkA6YETYTH216nKvSxid1nErx6QM/t33KGXRSlCD2Xs9KgYlsb2dff81d9nujFE+gGwc
+UBXDkLiy1uADjqzNB9u5vHMgi6B9JhMgBqNeyyLkqFg7x1ZwKlPkKK7r6Xk5dWUcQtpjZXyVbMd
+rM8DcI/62EkCz/u3QshsSMGuHwFaBOhfCZbwqIGr8mNjrHYiu5TlYXAFf+kBnTwtFaAQ3yR6fzq
K5ZRErzfTF7ctAnjOYzWhTMDkxUzTcia8TNqXAOsjXmYrMTjo3eOevxZAM8ZaWzyXOdxkttBwf0V
ClHMxK8bAjm52B9/CYL3fT4ddYVmdArzpUwAIoiUPTIS5ZjJ3f1HoII7F1Vckl2jH/KfFh04bf58
PKqNbULH0yyRD4e5KCI7KXkBJ7WhXBCe6olVBziSH60I4N6MhhmNErrx+18zqLmWr4wFvS2ew4a/
GF+udLLzmPT0lJgg/QjbphX71RtL6LFwjE052wzZurOnRYNoS/Dtd1EpdIvcPQrGSDu8B314Ux94
55AAirrXWjJv932MuEPNtC5cjpcSt2onA2j3RHcMXjpl1dbUB/zTErPt90R8oEI9k9qsA4+yZiJg
4dUtA4t2X35UHGbbBFItaz0xX2N8J+hQvIedaJPzLE3Xao2MvTAjc9zhcsfisrMeb/whkZQC4rIR
cTGyPqaJGhZMjNaJZ5nxwcgKYpeM3l9pLX/xYISAPfgwHcYLxNMBxcn9WTY1CFgf2FueiD5PaRZb
0fGVnM/9+9BygwS4ER/PjMQ0ZN+M5tJwPqTL6wGaAoM/BnkaIspMRtQaxxWiWuY5jf93G4o+ANbp
UZgNoSZFv9YdSm5bjzD/4LIHhG5XMGZP2kyQYgKofpKyn3eWUXhUVfkTg895Hsqdx+qI0jwrWQxD
waq+2f/hqs4sHmKHPJA90U/aHUDrn9wJVkl569G/8xZVfhZvBSpwSBAVKYeTWpf/a2Zxn3sxk/rx
IimCoimBEuNxsshcbezFnUtcukdSbQrNQqJiheOxuDf4gKmhMQoTFKwoxbsWYVHS2P6bFhiiWb0/
rA1hHTE2F2ZKbLNB7yScrOhyp96RIbNHRTHYUnb+bG3ZUe/5PFzqlNwvJJLJOGp8IS4d9SyP3g4G
+pPky/XDPfFa5D1Xo1/OhLqq9AwVHpqtEZPMSmLiJ7dqfujccJEjLvF1GLsMYzplAumqeoOWqNoY
jZeFvKnREfCpo1jpFo9tTduV3tGcdmE1A6YBxlQ0g8zG2YXiBMlgtP4s7sZuzLCTMIBqWRxVR331
SzHfkVRGq9pBqOAPMM/6jvQOE+K79F4fO+X3/A6i6SiCzKbcGv6DY0luXuUxbqRALyrgPwjID42F
m7UZbEDToE7I3k4yRHJGpF2tAAFzeyll4s7WWi43Pxkuz2Z9idmyzSBL4prT/rSqhnPzK1+KnjFo
Jv5K36oFL4WJZAykhUHSkZygADm20kMHDl9B+zTlfNNp27rQfFhzX/idmWWrAlN6JP5yUWyWD/Ll
4XulRXdeI5jfIgUz0+5DMWRzM0iZxJQh4B/KNtlc2YSCbJ6z+fhBOxRgzgtVlhkBMc8uilf4YYYK
rlxslhC55nqDT8mktRL0m/O0iEQm5EOplEnKpfcBxDqK1U7knmn+fS8cXA8BCedzv6hWsv2ozISF
ap+8qiVR35CuYX9KKm6kpfHKzERaALDHetm61qRlmsBPjGZOuSChDl8LUK6e12XaQS1hVwF6WkjP
wiLRegTbMJoO3odp8QqOyc45CY/rNgThGJbd3uSJM12qpupLAWi2Gs02SmCYN+8Yf2DkAbm8F8N1
FSnqunmlEcQOmJI/FGePb7k2+fesc1vCwlqlB4Y2WYLXLQA2bNk2eUADmSzm853EccppOX3ntEUo
0Y4iCeShRtMikfFQzCRGlbOADscIh4RZuq735BcrNdGL3lfZCzLyw+A86QE7sSjlJrmkBbg25sRS
VQl/S6PsY5bU3evO73PAkF2/6K4mJmmTcx9vr1cGRtX4WQdrZFhb+WuxEKSmO3YSoJWjlSrGfNrc
PK2MuGzZQW3XleervNNJJA84T8+7ABJ7+3Zh293PwS7RnMFCV+YS+TDlfutTXYsDKPLG+s/LCxbF
5lGehnuw3qFMdILwMOdPkKnM1B3P0evZSAGAlyxLeONaFbToR6Kr71UnqfSwd61slY6E5nLnPTRX
rjTUVgLo9NwkYxxmbbKFn/WZcDZvARFZoZmFHi61HIzYSRi4nKqN4teQN/edFdmdblBfBzLPMDh8
abcWDISSKxEGV6R5g9sg+22Se4z3iETakG+mz3J6couOXBhlyCMWVtt5WgF6V56HK1zJVymNwOJo
z9GcS6366wIxUJQpDY6TWiVw5uA9y2Gqxaz7/NEqy2dn8vNBIntYFRR2VxMPmKdHok0tBCQQf2/8
NU/40OTdnXT1eabK3Ig5qCbLNfIoMxmGXcxd+U9IXB2wt6Bcac/NIQVMSDjgvi1ZfBZPj1SsxICW
n0qmyfGPRKNvJeBLGqa9JPs+3Nvek8OAHdpWZW7WHKpx6/HQh4Hus3VZrYnQjMlNffNr+EDYTmUV
gN/vgniL3a0zDFp6Y526sPQJS3jU+rTeRXbpTp0n/BD9BNzB6ve0F58DW/sNpfVwWmh2nQ8OkUlP
vtxbZoytl6R23dEdVTLHtclLoePJenytCVcvnrcI5Ask4VBJT4SOhYtWIbOk3yrLi9vrQ4suibqO
jF6s+vlujgDWvMTuG6jX+kS+Yr67Rc/jJE2anjCvJwB9NPS9xgsFcGq7o5vmVqZfysIQwHQcX/Gi
26ntbIcc6HltOHB1lSjWnfZpxlf/l/QEnNkZArGgeXZBghj57X7hrlrHhR5tKEUux0D17fO2zcaG
RvpbzVuS7Q6uiMLwLn258JjWy4uoGssIpnOGs03blxkQHLpPS4xq7uH/mQMU3qaQ0O51Ta20FbFy
GqN2uOBfln4nNE6nrVDQhBZJ84XZWa8yAngC5Qlfe4WCIvftPDgi9r1ZCD0KJuJ5Kh61sbnisu6+
UcYkMVcxkXwKxoP6ada7ncbEQ5xOU3o8mtn89r/2EkMxb3DnEFP8NvvKOQuIZdJmxNeMPKGiLtdQ
n9LRAmPkXgrjT2elVEYSzBQ9yU2RJfTl7ldt1FPCZ8y7/78HAW61aoj0SRz2nZyeBJs2F/Pe4cH3
9Z/siqCnCLWhZh0GQkXKlhG+etVKSAJcWv1rJKXnHAn/1HK8xDxk4q/VO90755aiRZGDAUOeWey/
wbBfi9FTlgV2jQhWiMS19wV3bTmMnkTG6wFUKXsQV3vVDtGUf1RYMUF0hK5omsrlijMaSRLiQvYr
DP8Ql105B1Pj+17KKh2/9wi4ijsTIxmGFXii3NKtAo49NnpmpOiKsgzjmDRy27Eie62Oyn7xYZEt
7uNng3SdhqDm0+gkk1Eoyx8FD3xhK6v1FJqLb4kaHzwb7oh6+pN5hXiCBnFosJMLslkkP/4Hi2aV
zLnL9kse22o84xz0Wj+LREmPokI94i2zQZGh9sHYuTKVCJl8vK+gmtcHR6tC8htcOR1s3clHYstW
5Ra1To2W417UgrJdyXhAT+mhHVFAjQfLSV7wuEUXfl+/KG/ZNA3tGtOcxXXH7ca3VSowBsr1xTAo
Bj9lpvYUf6rlN95YSX6Xg7gM9ogJKOZ3OqUqg+eI+YEtDwpL8AwSLxVCSxp+/Rr5dJd4KLl2TFWg
LfKnt21kMksLrGElfBVyHoQJAM7kX7t0Oc39ioOzwAB7e44Cxw8of3w3wY7AcBpmlFXVIuqyU4Uy
l8S+Ogl9Z0khzq/Ws383n70wGbsNKlXBsXonPe6JcNEgBfmNlpOsz0pOz5Nz8n33P1qM1tlOneex
gRZ7R4L+H+epnG1tXrBP8lDIA4LvPug0qONa6WozxN7q4APmD/PkjQhDg0wLIcFqcNXGZRQw+rBF
VvEBB+UVOvdquACApqKooewWAaAxuRAxIBS2CLhH9o9dNxgcFx1+Tge/dEjWLeWYgatR9CRDKXjT
V8faHLEF3paBeAA7A2jobtzclEFURbJ/4Xs686m7pguW5+KhI84VaYbwdWP5u8p8sZ7vK08NQWxZ
Lde1TJy798k5V++CfhQEhRWSh+wfpyDcOBiWF/Lqz+/EATstHWMdWz34po77BQ2Mq3sMN2rDQoDQ
23w5MnlA9Dlzxs9I3cJ36Jht5k3Mk77UVXrLj45oDOKmGJHfHZB8pY5bh+l9/Ze+kGmI9PVymfqC
/ZcXjYx/F7S4ydP+E6ANwbXx1Q6QAfO/holuIlsR/0axfaYRm1A7GxowFdWBDF0Sj8/0Nn+7qwFx
Kz/Nm5mrfxE8qY18Ar3FfNaFPr/iD/wiNAGSVCdgDxX4l9Bjc+/001CJ60x8vU7d7rM67giEPolf
UWIZDMtahY5UdOdkkodyX+cTdJKa9K8BbkAnz+LGxS9hbsHyN9ncaZl4yi8p6HGhQZWWJ79+RpP/
fTjBWZLU5pP6j7nmyA+twPCaSKOKjsZPaxyeXd6Z7tcEo25xnQRG1LnyTLZ+EStXXaHnmChMKMy3
mQqPkWJn4wwl7X/6eO1vKvSfBxuykbdGXo7ggAgvAMqFLfK8URCmKgVWN4GOxuUcGomqqNVttcDr
vqs+SvaX3I4JCT9VmkNyuo1lMUsua9cDarP1kiScWiSpubpCUy+Bm3s5q+RJZgtrL52U7Cl0lA6M
w5GBBBHorMlZpnN0U81obl0IGVxrQTcaxPWmoFCKUtr1ioMuDDwxkLJGDVvgNvrbro6GfxYw7/QW
RLKxhxxHr/BO7JhRquU2wXTk5oXbEwcahenJ14QrLGKsH0N44piZwE3Y57R7je2eUVc8GU1nb/MF
4we3fC7AIBC6Rqz0guinan7BGMcWt/Cykv5N1onygiABWHdBEwFuP12ML40FA0kfcsyx14RDUD5X
bjg76FmOwh3lar6ql4qO6ZxJwmygLHa6qhb9OgP1eieTBzqVllxbDLY1q7IHIuJ/ltQSXkKtruIT
gobIn5wqK3abV+L7rowQXkkVmVBlB0Yq4ffODrlrmWRy3qLbi+t2n9zYWY0DSCPFcaMhOQS+jz+0
tGgtKcYtFFbwKrignjXZ6FNOzw4aWo6zLMyICWnzsGjMUjdGHonRtJv3ySt04727VuVwO0qlociL
2AHOLgSib+bvMDI3nl/YP266AuadDoAjg7FI680qqFa6/SShBKutShz905zrfLP2OfgGJz20vQih
ZHF17kbVH42rGuAx5I5+vbWW5Mu6QxeABfUY76KdZ7c3lFo3OhM+mRuvOw9Dt0p+TsaxFSU/jPES
q5cDndkGKtTLhWKQVFl2i3BjMYsXVmyIu7AMV3VJ1Sc+e6mjERQZ+WBLKHPJs347Z7oJXI+Z2GIc
WBnP0f1o8ngUriVMtKwuK/ZNcuV7wj1PdXJq9IHFfE43N6fRp4FMHYPkCLWwDOjP5AW8hCrKMjeS
XUe9LRauNJBRK7OKx9S/mtbVHa1HhVO5IieiCvA4FlagHOhdqFghvUyoIRgsi9nEWBijAHTPyjla
1pOhJOhAxXQLcGPiwLJ6J3FzTzzelcCTXhcAGAW6bmtn/2VvdRGGpLXvPW1CZW7bYgmhPmO2Y9hl
WS73qly9HgnCqop0DLwIu/ES6jME2mBUn8Ot03g5wd4g9LnWRUKfG9cre7SifyosS7xrNzWm/lj3
M2n1pXFVaheVKUJpa4FFnJ5GGrqwYRCvC2sHzRAgNVjzss6iYatzgDfFxer+Ock+L/zY/MGiUY5c
SGqliskKGKJDa/aM0aJDlaPePpbJnLM7v93NVW8+hHJfyVkZyJHEBzVNO1fzLusiQA+N9KAa1C45
nqXxo30CA2EfLJEgyn6gALjqurywMVNrqgsCQZdSJhMT56zVWrzfYtBO2TL7AOXJegqfDErwYIWr
hn+G54OthgoZrmvaECJmX6sueI28i9MVMBSmzW2tUXEimqPO9Ahwuga2ToqHbyL7YtVY1x3oulVM
Z9UxMFr3kVxfbqRP97/ApMBFIip22uJP1HckLQrBjKerNQ13bWJKyBMEMhzUtpekesVu6h/hA55F
5+HxbMNLpZZuWPPiyrZ4GaGXiHWxSKDtbpQvEbbSNuPIBMmEqRqxM89Zlxh+KoJlsfw1LdXGiaaC
g54pSq+qBG1NZctlFAV91H498gFPkHpnu0kJrbfuIZa4Kpt3yZTxzP+VQqQ3bvgM2HkgTn/nuJ+6
0+ONhWsO4COiUqGis28csD5iqS83JUGyaIyVEoQQJwf31iqRjOEvQAV68TL2RV3VZffBVtmtC2KR
pIIBBepkJ4weTWyYyIidyNPdmqwyN4tZfsNud3rAt0KUNIVSXt7TtfRk5N0BNvGQD3SktB7LKgOz
GywzHjIbSQ1vIEtvi2DJ5YtTrAlnCT+2wRgX09K+pFFVP35btCUTUa+0aac/tvAWmpPj+BI3fpR6
f45RFrrAZ1b9rJcwTjFWTBOWlJ09yKKI4/MCPbelhi7+qiLLh7mMURsgT7RY0UzuFQnFUxtve01v
aDKM+7oWyUQGmaJ7pLpmzFnucfE3dv8Ckx97OCH5n/ILCCgbgSAy5AYC7a0oASctM+55uu3Zf75j
nJ4akGbTgOXGB6oYKfd2HpA3fJQInTfS5lFReFb5rYTPGarA6aBk6pl2WNrrDxrhagastbv3IMYA
/c+pkr87NTvYuxlBIwePNC+cVjyYDsZjzKnppLS5qbsQpGxSU3j7nqDStfu71QmPGSPOFrZLQEKK
RqnK5UGNaBigU2xX5JuC3LS3ir2YQeoBPV9SrfgpNdxkuRBd8ImHeldQlRNNQR79RwCzTRxrcp4u
dhpVEh5cReC6Hc7+AkgQC6OUfrRvL4B6ZvQHCuJgiKZvH/yAMGAYHeIogzLaelpGddDiUZQIIEnc
nwvRNGOoYk5cxExI9q89M8BzrAlelwgXrjLcz8ZOBrS9tWKX4GnS5RmeAdK557/Bzt9azU7IkWeI
Oa/womAhwSyxVtEm7o6DJcv/ngv148b9xn5JEc0Dquegyr6fGgu0rHo49Hes5aYPC7hOq+WLVJLl
n0/CBcqhLBFI5Z0XxF8RC+71wVQwDDWYbtt0u9DIGtDGC2sMn42+J6ZyKGQth5TUDXzZMTVBKD7Z
VMc67pFR7giJ7QyJc+6zG0h16i6Iva9n1EyPLzlGrEQacxr1ULRivxMm6G7YH6VgO6TbC+SCVfeF
UZZ9ghxWc7NiqR3QUTXF6TtLrfHrO8gTTpCxyW4CVsq73+nvN6M/ehf8cnecTT6s8yCHmD1KJrs+
uQPjkUpq2qvADSGpKkywHiDvSdAJ2AlGCdcFknN4lBzpgD9GNMNqHt5ZrBWfMInACG1jEUpZUd2n
lv4BZUbkp4FXSWTYoJFoHKqLxkOSdeTM6VyhdOxh4kbv63634e+kZ+C17MU3sZnIwKPneGXtW55Q
T2MBwKPDsTEQyq6lfLYv8fxGiOKjuKxvJT4W/KmZwjldp1DF+rHn/XeABVPI+exb+2z8VyGiSzxF
TkN4bf3kD4vhOIGYqEnhM2Tuk6kC4pg8gpw1txsBJV/DLckTvGujASnLuzqIT0P4u0m/8FUGueVa
k0CSYaAKzs7R30BBgYBbqVduux6y2OryYVi0qLT8Xd4+WlJFlvWxJU1eEgQfeNGEFFHqot+Ao4pw
8thGUU+ZcmUFJKPYf0QhqCWlfadySkKVHuBoNYIzdTHJ9K67JqYKffuPUboQsHZnbcOyQqkfFtpF
cXfbZS2+eZQxuYRHrRX9jY8PSiGySw6jUVKVXPgsxDBZPzTO35FujxGqbkMk2jdQ+u/pYqZQYLGK
Nuryo9gEZiwNfGT6LI5f+4EJXRv7iRVBFqP6VTm1bVYO4Z9m9yi38XPx3PIf4m7CRSdV4Thm3iMF
+Qa4zpCFEH+snrCzmg2k+Xtqp+s4OIuJHkhAB0Y12FwsKW+MmqtNHV6izXoyjzTSd4qOgcNxQIQl
idpu9spq2Eax/Kr/uaeHP2+D+j5DXr0T28l/alcYjkioLRCUtcRKMREvkFkuIyaZ2KRRQlnO9WlG
fHx1eZvZXjfZedAPaPMT1Z5lERWIx0BxJEd31NPtt62jMBolEj6du+WGT+XKaLw4sv6O7/F6ld/p
1xn1dcuYT46MWKhBfEVlEJRaUhaBRKCUKkmKrU6JVB0P08Exrm+I76UYzqCuqux4TSSziYqmtAQb
1ilFz9sKGMX1tGiE8JzsO6Z8XV+U9Lc1QHJ4IBZH+tT0Z8lOSP1M9oAGh87AxBi9nuaFYMlqQBob
CWSVyv+vWIkTcvXKo0i3H7oh4Wz1YNGqN4hNZ8Nl4cZfosvkInOnk4VG+pGmi/UTzxnRgjiHlMzc
YYQhMYSxdqNOPybzWkKLvA2g3RPECsNHgB6K4sxpSFSTRAdJl68WtxAiZxp/1EhIACB7TXSKFy5t
ZDCjKmqfTVnyypiJdGnpfN48j+sou9tX4kPiv9Ih9DMJRiHUH8qe1MTbzSbY9nay9JD2K6dC9oVg
mwZyK7OarDQK2bSkosuORE/4JKS09O6jx0nEwWr96Lj/XvISgWcDz9TWhakeT0uwKeKglXw3/H6F
cWZTug1ip842iTQr+jd8bysyze/gsUeOcOC3iil9WMFD/BXINJInVhtnJZKPwOZjXVyTnBKY3++y
LqP9HgKyiSfkgWWswRHQIeL7T6ad4KwBXhp7FU9khe52j7/+vPeACWyXQ0RtIvh/nlYlK95dgrM/
oyjpUhzYjcsRrxa0mtRbKYwK+IAtO6rzoHKB64Hc76nC62Lo3JB0LEvpwqiP0YMRcAMILeMcuBkS
eGjulXg3X4Hw1jVOAYfKeD0NUB399przyIr/rhJf3pPE3P7FriM242TD+SJivQWyhj2ZstFxVfQx
TeObzTPZeb2bKFi2kkqAbDxJPLlVKKgd1mK8c5JDwxIUNo919FcqmWrtAOE+AlqFks0H6baKBXOX
dL3K+3YQvysPHId+09pbT7pu+4wVzfJKLgYBnv2qyMHgygvu3f3ckO/Z8+hu5DgFdGFauVIGZZzv
X3iNnAIImeV4GAtaN3kk1BwFnvapwNt/qZOlIuJ054GPM4F2Eqlo7JdQSHkNjF6e3EYhIRak2XhY
XQlDSq9x/GmDcxmMqPS7Ylw1qk0gqREPC8lO9VldXQtLXKSsr5KQs5T/L0/CcB5OXA839pb9Y1MM
iIZkEEWisebA1ATQ/XkAo/c2DjvLjTNqX92VlOCnm5/kc0aKxLtmSPF8W7FzNzmHrRL/LAYoNiWB
tK1Tyvj1fm/SIyuckLGdFz9QPiW9h6BcVJR/b4PuEyhBqYhCmNnDwQSQ8iWfUi0OqXt9wCywaXtE
j02Bl0+p34dUnbUWAOGQQsi9nKUX3AtbQhBRd12bykGg0Hp5ATePJoKyS1v04shfoXBFSLxgHfsf
Twek75TCkddosR38KCGT+g6WOYOPg6QPXP2DdWOULPLewR2a2gwAjM57RPA2tYNRDSCnJ5VITjMc
D9t4R4tbVnEVFEe3xHaMYHJda/bcziL2nPDVtJIdSx5xDVRKTaLTtZWiPak1kNfUBgRlbmWVyjar
BgpjO8plcIyBML/bP1LXMzUYqH6LqFUxVCqMFNLM4smgeJvUuBnFNeM9OXZd4rINGN1F0bMgDXb/
PtxCnGR7IqxhozA2Qikad+dtyMLmOTIDcKY3bY8gv/90hg8xPSttOcEXk8tt9yT94H7X663YUB2r
B420I5UWbAdqECBvaeKynQ50O1JXzwTHFp7SPYhELp/gPFUQmgBGbJSfi7XUnRzHc8kg3+YwLml9
GjK5gTwB3IFM9Hy5wBAOyRpX4/NO4oYiya8QgFWUGGaeT4cU9cWmaHpEWs1nkcYsKVOZD3sM6leM
DFWNItuBgPfgnW7YkUJO7+5HkqvEY/AN4azC+MBpxzRMunCmG0ufMju7umFxz8Wg6oG8s/ETds8n
Fuu5M+iAEefcb7bdgGc27m6AjyVmdIIaqWGAn0xV9wJ4g/nrpyphlY9YIIc3Fwks7ZwvHwrHFyaH
6irn5+wR2hPQrdsDdNrAQpXsG/Xv8x1svPP0xUclkQEl05sRN85hrLtdCOt5yyHwfYQB1lbT5l0Q
aVbtBM8QIulOKioJxYmkhDz/YJ4SwfdKr2ygfqdMoplf+p8ZlF8rtDkddDvuL1EgEnnVs0KsFwoM
ecE+jPYgN1w25xdt8/65JnbQGdcPNaZhq8kezJDPpj9+VDbC5ND8SPJB46vhu1zIkGBHDfbaWs5D
xGnSXvICTOdQBywq3wXPp6YVga8BYnQgdzRaomueNXYiiSvQuIyPTDPeHCOgKbkhfkVjuk3myizL
vS+cGlwzsvnbTJxM0YGCm9GHHbW0/bXJ1FarSUrqpVXe+WZaVCgQXlEgcBof8E8f/4xzW+3UvwsV
Yul3jpGvfmD10GRmgoFf93PU+2yqOAOiDre8/qZxFE2U9fnbxnKon9C/pNjioIdKp/yJUi99Qpnk
v3CSFqN4AEGJp7pNIKjGgZqO2R2CS3asiVxB+wWhjwH65MleMnrH0b/IQ1V5R/AEg/x+au3tP+bf
cKEZ2qnrgEB9LlyYzMBHcA45jHENcnVK24qgC9YG269omX8q4xTb2xbUhJJeJkgIeXxblhlDrEK5
dOBG3nqBuhk+HuMrknYnZQRJs+3zEQCUFZe/n9EyJGCmaPs1b7aHz6abQEeUmgijaXeO4YTm58VB
fEqYOicne5nPU8eUMFg/1AweFj682kkCTE2KKiYyy+C/Fm22/QNDIrF0VGQw2OsLVqGQmSbEjHDW
a0BOoVjtchnYTwLQifSBY3kqrm7emY6z+n6HurYjx5EvOQjuNwZDGwYWcx79LgCLjubIbW+8/Uk/
au09HtCDTgFvBkfCyaeVw/GKba34Qmi87V3ZxFKwye8KPOFqJyWsvmT8nYsGMEHXdm0yKB/k88se
mo/oyf1lpW+Dee2K2KTxASJj4ftuzyPeL8Ve35dWxFPgl7knNU1HaW7/W5dQQ4V4zn0akoSAQeY4
BAjwhg1Baj2YXIgrsFPanFfaJaOZgJWWwjMl3bdJiCJpfhCHgDs+Zu1rYgGl9PnNgfHu+iUT/eeN
po2N/ondN9XWUMFaQ/XL/za3eVvvzVHM+5W78WQyLu+5KAOo5gbIphOQ+wcL6LsewU4IdLuU0/9E
x+5PC3e7z8Vz6wk0F0zGR5Ysoz00Fa72hOBbCS+hmBtcdCVxCkGifj12vZbM2jvAlHCC53SpwiR8
smZfPTTU9m/2et94BptOPAY+jTJXmK8YzMjZK4DrNYiQhMs8Je2Qh0FtBn4321HrnInPelKomdE9
Ir/sf5Zn+s6brBXbaQgFP38E7+oVPDkxlSQ1rFKUUXw6pvGJ4QvE0jV8OY4Q9v40gwG/4UkSQuoq
6nD0xM7KwyKkEg67DiVgHA0kbfZwu/0F1+APdYxXJP9ZJCA7keyz0NJPLz15KUJkKSvPLXkmM63s
vgFDM0HchSvgW8TOcUCgjfz8vLpW/rKYKdzolIBCaoLliohNyk74/KgmMPVMfh1ZKPCy/O8tNIJw
dSzLA130IDtTOcMzwV7/xcpnnLtObkHDMpWacUDq6Rq8tssWYz19UV4j9bD9iKRNj5bWq+2dnnOP
sjT6u0u53NusEYYRWoZlEWc2Xk/a0721vp9yb2EEM+LODHxKdOCcD5DtsNAsy4mIDeZAYpnNblq0
GL6i3FMXHf73PASlU4A8Fo675rrwgWQOlrUM6/t5QjtlGeeTF9/D+SkuSZ56hLpQnb+eL8CaG4sV
ZBG6uiVvTMUuNFnY0kx6deBxcmySsAXKLy9QmdScKw9fjDanmCrvzgA/7udLCnmWWmShKQ+HUlYV
3LiYjNGF+WgC8HDKCDB+CNuLx14ZKP9F2Rg2RTaO9eHRNKdtn1OKFX2fpbsicHUjnVzhZZRAbbHf
RKqjxMCx0ZwA/stlG0lcFD260DaOcBjkEqJmcdTxg7ZfthlwO2WByWfq/tl/3n4FLi1EEtgsbW9E
REzZRaDLQkA3ox+e91gU38iy7rPEGkNJ0Pl+p+Xtx58LFHzKHWi9MM7gfGwPQz45gtIb3TEwFjX3
3JWa3oF5+KFUe8mncvb0t+uvUyVwNsiZ01BoIoJuQnGuNGXfOTeuOo7DB52YnldzkXzNsUyLYReC
XCaYtzJ4sTxLDfKSUg5inpSjJU36Q2Txn7ghp496HL1Pj64RJPqT7GBat6BaWdhZNadlF4JRpUjN
vwolO2XHBPpIt09tFOpqXY4ZvbXOKnwXIDu6bw8VPxp7NinEzevqvi5mPoi5vqnWVwSfMg6vm3S5
DMcCCvgZJ6KHQxP9flgy9P9zp3ICza3IX60WOsQsfnQquBJAb0W7ZtVmH+Gafe0Um3tfE4pVgq72
dOXIyzg/suvUIoQtxYq6agvf3hbmuWBcxsQKl1w6F0xSPkN1oqeIeBjz7xQIxt5/dHilCSHOiJGI
oZbdqPklR3x9vLlGvrUTIXkCrKeLXH5KVzc/wzxbE5lofG5pXIHdl5U4UiZY5AbNgMs9evhUrIVS
B+fYEEayOUzFLcKMu2GkXqepNJmMAoMwyI8Bw7ZA8iRxEq8UWypalAxIZqJPGpZu1QlloNeA3Tj+
zXje9fk0UueQ3LFNfKnEwGcuZCY9W7SYGdCWCTTLNcVFpjIBsmHRKLO254zaxITJaxJ7JTFrpH2O
oXU/cY9HtVzyWWEw7gRRzuchJpBn5Wp+QVdWyZG8wUIIITXaJwNgrNRuJzpWDMupCIWL/eUlHQLZ
O7CKHqxKkqxVkP29qGEJ1dTJ0T/tTpTZekuSVqYiIMnwBxM5Mj6LMQPpXpGL8XtmNI9KtAQz8rdD
g/vuv4shbdjlvQeuaQWeSaNrZuCuU0U/xCL8NL/GpXBHlkpRRd654TYh6cV80sAiQtp/12xJD2nB
Xk/jwxjsHeFJqFt35lqaMzRwLcStxLA+53+pYfTAHYqUjx4xSNaJuF71Mzgp4YboPCE22+qlflVO
jaMtem0xirlVzKrTfff2sBEScLJCUfD0RhwFXLEFupM5Z2kPw4wIzzsWth7gFqYpIAavmO3ngIEL
sgc/RkbtTVvip+pd/VoGk7iSNGF64cvSoA0zc6Se2f/59xYCcEB6zlzU9WSrsQ6Gfi/p2SyFZR+5
Vrz4FzciHJVB+loQsxbWYXS8hDL/g6YtfHAI5E5RDZDMmwnIR9FtwIlUPhhFWFhTUmqozMNfCQ6I
XLzRlfrzoL924sKMrsSf3s7IaaSzGLA2Fr9FuB6V+Er4oFB9zsUeFrKAQIuGnqxjbxzmeg3lG1sG
kDU7rbdvGkHbbNWc1iBuqztdAmsM7eGA2xfWTCe/h0E4HaouFCrOz0QwhYPe8JPxdameB3+k1dRZ
Hegg3LpTLbKAj00hqgvxQ4Z2zhjpYAJAaOcCdUEd27dzrVmSUnMSGVlFlWFrY7hZyd2kj/b19Dtl
jGjIPqGBJh7410nlY23vyh/S4t+GdIOP79dMtCxGPd3INUki/NAX0QxsQaMT1cVVdGG2KNr8UNNT
VW8dBTB5g1fDxpzSAjgyMic/nlSrqIOyM14w65DyvDqJDBUvPqMGRRUtEAmyCkjmt8YZjtSUFOKX
wzCma61ExhvRzWlKwFXGOL7O+tgiZk0hCyhkYl66XV0WssXCcJZBhf+g1byMywyX0BBHS5vHfyqg
UhJPYLTD27Y+pXNsNlhbmzu8JZFm8CnnyDD0geOhkAOW1z6kQzEpfan7S/tXzM4jKWuAOK1EdYuR
GXZfKmW+JLfB7HsBGR4JVP4WKDDT/gzJvgqYFxd2odMsYjBXbMJYvvRWXQYOnnqCiEFogs+nKWW1
RhV0b2zVrH9LbA3ogOLGRtBXG6wQyNgks48fqFc2rIXZ+ccm0P16uqW55omFQebCKx3KKlLyJQ+/
xFxQybIDQ1favjHRB8Kt6d5rrgIZFbzFf4FBLl3kDZ5l1qVKcnRJuJxxWipgUmZCPw9c0YHJHNjU
IzzW6qUKelhYroM/Pk3d32I2hkgbtPYBeqXJ3ndjFPZkl3e3zDvEOG1ZNX3Ps8TLgE9qU+HhVQpM
cWyu+IP+iePwgC/+jbW+qLaHsCGoVvF3u2AfZOvCD9+OwJsqR20FdenDYMXKFvxaTYuIVfD/+EgK
/2xVeLHcJf036IKR1PuuTIGDhj4YA2+OdskKx89goalS0I7uwajRqUDlr1Mc1hWt+FlCHry+WAlN
aqAuOuvxvxcEY2PlFp4Pr5EbMgPvAO34fbapCOQw+WsQMwU7WX1vqaRgaef9lqEW1g429ekDHZwX
45jZu5/lbOkWbDRKMn3nf6wyFjNRpl9e0GllJuz54lxb7MaMZSFUoXy71M5xUQCJlSy3X5Ix9RY9
ZOqvLYqQOLVQFYoRIQY5aN50QjFE+qntVJEBEMR5GaF8Ymu788hXiaeaNvQfu9wxdGwykh5g/Zto
02xnzOUGCEsHP9ZGespGXlPm8TdjUKeVhN4U0q0G8V8C7vpz6Q4qNEca7SZfON5E+6B77jMt34tL
tm/y9wCscH6TckvJMe0xoIL2TMvMNMe/TyVN6ipV+h2y0/E8MVU0cYF9IZccGcL6fiAx8MvPQ5eb
8HMcEtJBX1Sa+cnhMBtsLGMbFhgawlG7coxWs0mvzNvtUmPsF+9o88uuINMfsMltVwouXoRU1DmG
WZ15NTp6tQ/ygwtX7yNN+Doh9qhjg3LBMdGtlgDQuVh02fNhjno9gGVL5OJhxyJ+s5VkeNJv2MBD
q7DO+JsX12GYrcYOyfqkbwWBFQtGbnrmW7JTB0oTLAsL30JYpxQ1EzJLHm5MdI1yhsp4S0JuaTdV
jW4yafxoFPE6Hsml8VbwD0Lgx5jkTraye7mhCtzsy+nGtPy2SwYF/LUETnaA1iVyIEJGuqtoyWI2
njEmUzdmlRq/wbzUHfDtahtttnWm/n00nMQ1mFa9hqyJ904GZnNxOGKHWA6LEVO6j1KTDtvkxMg+
YYeGTb1KVT49/rgOnl0ydhFCxcrNE2jEYTcL0TvXFC6ni8elHti8z6ndC5x0Xml9b+CkTGP1j+GK
9SxjP/T0My1V/HFm4h4w/WKGTU4Ejq9KCmEOOmMlHuF3BQJTBUyCblQbcb2FzRkSa70ffyIuBOqS
xPBYQUBUGArQ5WAdh/dMtY8AtkWcoRa/sV9vXCemxZRh5VuimBrKy66reQQInOqxjmaXpxjeYOYt
84e8sIaBPwKWA6wA9FuSd2BUvRV9d1NqBLAvvPyL0K/xW+59UWjW63jT5/ddJ//LJnu4aBiViKmG
b10TtMsQiNpdjjVySJ/uuNGmlbJ+n4wVyyKnsRKzugmUec911QYXcJhGrgHIq/dQChfyg0gsURdy
MvwhKikSFZyq3T+IvT/Gemf7yPixhfDQw38soDaHK3/Q6rNTuXsNhqw2U4wQZhlyc0F7Zu8lETH5
A7qWD6OKMKaS4WOoGaev7obmsSrhS1i/XFFz/zJ+L+N4D1DdTAQe4poP2oXMkWDcllIt4w7sNv0Q
CIZZYGVH8J8INMEDOG/udrRgE3YUtDBKFhafCJBckT7Fi1XLg/8Z/JkgejuFTRpwDhx1UuzWctHL
d+Ys+iCdINIifTvJ34hNzMzXimqDAgmf4SrOIMmLlR/7qDNQBeqVtRiM9KdvO1ZahvzIp96QiGBw
Lf3T/xMgQ92Gr6Vevux06/WEL0TYVH9nQN1yNR4yQJ+Y5giFDcil+S4L9G53sZnyxzziVs4V36YD
MB3v/AtIFXpS0acYR4H3JAOH5+Jm/3yEMyI46yuLHE4IHoq/Jev/+bt0pRKb0gwJt4e9F0hGh54s
RclEQBTmRenV+sisOdyGQQ/h97BQIkGGpmEgKDBVh2mHtuIC+6fu4OMpjvw6Lp9z8K2ugQ5niW0r
BJtD5syTmcgDMwrQQgfOStkRZpzhO2eSNHXish+uyI+D1XUuONyTRqqG47oIRfyBliW9K+RlrrCs
HenUm5fegqziKGn+BYwMLsiCqip+9mEWGVPBY5Q3dQ0Q3TyvqpkKIoIBCh23y8cFHBHvPS+vhhqF
GD7JuTWuq9r4+VGK/C3ZnHYYt335MD8A/mc2NHBwlk0T3oJkTzRbtrnQB0ht63mzwvzIaobwD0H2
WagybGLJmMj9X91Yn1gcNo3nhwwPKxJIpHYq8IMc1K4CRohrwiggpkuUtlqljiKkzOqOU9G9NIk/
Mb4Gy6G3WNT5envNeB34xzp/wn4+x+FWzK3tUvuw/+cXP9Yx4QiLUyMMMHQhvrVZYqowWE/05uke
GMQvl1Re4Og9OKruZqO3oLAmlc63e1NcTT2syaZ6fF+au49AF4sClwGgLUUCJ6ozj2WRnYastRyz
aLahB/45NmJ/iKSwcy8LYXx//tiMutTOBlZJWEVE/TVKw/hNd+EskR2Q4S6kmhsRzHrOTkjyafNF
DtdQnDMy2Kqm0b/rNcpXxK6T8nW7Bz/JPvIaRW11IeoN36Wrw8ktvjxceIlmUQGyf7BEVCIEJ7gB
Ydxx9N9ZZhBiyxGo7DgK8+oNS5Jx5mBKjcVFtFc4f6znX1hg2tUubmYrNvzfjOV3oAcV4qeoo+Ga
oRKBkog6gatKEhkg0D1SgR18MqT+KdL+Sut2AxwRhcuUd75O0vR/j/BfWYH7iE4dNGW7kjzecWUS
Kg+Q00y/swoG7siHJ/W0VLK/XOraeyz/NieJLepc9eFxu9B72ln4m1VFnS+LAHd34hYEWwN0saba
/m/oWKL8/GuAjjAjnsFv2e3aRsj79xqHr9AWG+IfoF9h9QtqyZxY3WVNxXnqeu8a/KQMeP6ipnCS
zFPXgEryr4zFssGePON0qQPc3V9aKn72oLgUlokBW+gnClIodGGb8bOzwmBPXMp53aIzqqBWrLVl
VXQAqMj7AY0RCsAUqbj5t3ImGt4Cqt0Rdpt8pKs4FL1inVtSsC6kgFoeJCa6vGkFurk6/OnnwUgE
KD3j9nKp+8lBjmc6V8VnqcUN6KUkXdlLTmM3pvAAebq9HH2lpMGEpLp4iJTvZwDd+Oz5Ef1VLwmQ
W5w3INj8844ScGv5orcYc2KtCxPJm888dIU3EgeEWP/Vd3Md9ut12x0YtmnDm23fN2cbB/OjzXTy
JTN/B4SR3RvXeE41ZDDUOYXr9cqaFBcKM2SOvmmXPcpue2WhoOGteyrah+vDTN9bZvna3MKMfcEo
guoEYbCyK1zute/36Jkx/FR2IOoVJLxX0dPxpaFbdq1qGuPbjSXBvoEt2m+/qikF4IkNmcuDfTb7
bJm4NEIHhPEt0jsw1peBulTdHKIo5asbERqk8gdfyTOq5v062uUYg/1TV0xFuzBn1sHAU01wXwyx
UvZc1LT97RZCXZgLYcf2/OmrBGU993RV14KD/afGPxxA6p6/Ny2MBHvRmt4l8hsY23FQbQPALP9+
gFIqaeX11Z1p3g8TmNADHN4DNzJr5S5waAOq5LPSf5WjDkZfV59X7KxGbz+Eapku23kIJAFTDQdj
GLONFBnn/gmZQwmpT7WQ5k2oXoCASBwjeV5bhW9P7CVSebidRG7SvpOhNHe882FIG5+661JeCIWm
taHQYoOai8JMHIouWjKHdKtYF1uUxaCw8EXGxDgkiUfP2U7+/X63ybcx5VmISBbLs9jlXkSNRIRw
jfnMxtK1kebfUdWm5faKyccX+fvphYw0YAkXfRS2WhrGEmzAw44t6Ovkdr5oBE+YSfxluw99mOJ6
R6vo1BcJBd3bTOAc44zpQ1tF3UQbAMhpBFZdjrfg84wyqKfcmukNgRzTIv0uyTqvsgihC/SrzaOY
SDB7SyAdI5m/f7gOrqzKps/ae4hpUclaZ3tGr4ar88vkQvJVrvAvVw3pGD5ozHtBTAeOWntfR0Te
8Xe1t8sv2AftlEo3YgIyAVh9igzsyFcgYJvHmbMjw28ji6ntDTfIrGCExadKNXAp59ueTjo9a6T9
85MGJXAy/9SqGLLwfU39PwSZJX3sU6y9Yb/yEfooENUxZAYsMgs2l91fU7K2drjmCck2K/Q3wC7T
/Fq9N6BDZeGIyK1KHqZDMgK4Oles9luRmHUBuiXR5FUlm6LQNhbuSnUFuV/O7xG0ZpiP7RyWBFpC
S6z4JMGokns3biXZ4fNZUxvxkV/wn14QFnaLFQg6uKZY2VfBBRj8QsR3gCglwHYJjD/BF0Xwg5FR
wKGVkei+MHYJwbtMYKj0BidpIccGCwoY+3puKsBRcL7G2jlAOGiHBmDecDleIVECcxLsz2OD8qjd
vTNrJ1KF1k7Sd3Ta0Gwm6NxnjCH5nK4KMmcvPGNHyc8j12Ek9V4oDtXed4ZVAvL8lHgI0ylpStxb
AEmV4reer5QCZ72wE5qhOXUmEdTyEDUdRa7NlWDX9JcTnYSm/cDSO99YRVK4DxjNbuHQdUXhxnZS
D07qwmG+vfuxd6/lwPHNHc3xRCTHVXUNbT4JleL1h/Yr3eh8+AqErsra3YPWERWzXsFVNX5FNhCA
ByoNqMQ7w5E5n9ARQ3R/zm6uoh/tCg1FVIPmdJ5nqxrwZJYhFwDxfqaPHvCRPKuAzHjIy1xS5oRU
tgdNawETnQQec9jkCVOEL71ScR+7FDXWnfKNzSz41w78ibXR9P/mM5KkFz5DiMMJZ9bci03w/dfj
gmXlo57GZ5z+OYuf22BbvRgT+HANVo2icBCR9rhcr2GBT0JLqdrOhc8IgBDYo5mnghTNKkSOVQVG
9WJZqZVz8eMsxI6pa2ylGJcIExX8AT4x1UPwSheZx5W3YxKYUFRNFebo8kZ6P2h8gjEatoRcA/II
MFQIhuzCa8nagLNEhTsxxANUHs3eRQVHRGJ9Ppa2YdTge38CNI8oukqtlMaAr7wpcri1HITKqv0N
8jiDOd7SiT+8YirNWV5Fe//NoeQNDR67ZKheubme32DIwYljJ16gvmWdPefU4ATRjViSUjkr4jAO
rvI2Bn6gq/cdvTS2akJTFKRQsXJ+GYt9Ojp2Eznp5rQVxlhiv439ho1qyTIJXx5MHN9lwfzBgOHW
VWBeehijmuoGyjDxl21u8A2Mxli6qZM9QIqDo7R/JUpLwdhuVaLxYfywuaNg9Yk1Vfzx4BnyiEt+
GcRpNFLE7idsjcMZBYH6HF454ScxVhVaKw6xgIds8giwtDEzPP17uK8xrDoJEceylkdXVcFB39iF
P5Y9Ekd3XrkEdr4CA7528IxWPvnoA03rGLJgwf2+Ha72u/PTSixscpJxg+aYTgn1CJwwRqTx5RhD
WKiP/gD+GZOUU7k5RXttlKy3KXbtjVgtPrkN94HaZP8zuhxbZC7HiCAF1fboyrsZ0uvLRZV1ma1m
DSFGEoduXXHnm/OC8ym+Ev2zt2zN1/wtUQNUUBq36N80BdNFfDcSPEudfPNoq3ayLjLQeU6utmgR
+GCzXSrNZe9umSyxp0lJbLTPLhw1RrNG+OtTTHw0iyPD6RjynRafyY4U0Qr2u+qTvtqoN/cMh7gr
lT8ScyYJCLfzDyslFtGeXPWOG0rCPdy5X5fu5t18+4ugvEhYlJA2R93ZJ/bO5mEbuDl1mVTbu0rm
SaiaZa6IKgQbPUFABz4NXH79qrBjYtEyzOQHTaqmxfv3rSqKh4d0eXw7Wfdy7vtf1vyrD4CMaWaU
gJ46lTJED0tIQyN/DUSy11uFrgZoRqYOjTuY02X5cgdDgcyhNkHdd6fiqC1OFhCjj4HZdDYEtXqx
uULGzQSgg6YCFOWTOOsbE4JwY2QdIuGXVMxsdEQ7QHFhrgDXm+tpZMQ3dYZtoW4gG7b0g3fN04jk
jhQH7xO5+Y2zLHMPxn6tpMZEWZMze2xVNApbbjRPY2OarmSyO1JtiF9Z7CzPs1IHDasLPOiwYNqp
Tgxj8TL1shBTd+5iwq0xkJ21uyonR+KwFEdQtjycn0PsAdjchlNa3B5T2TeX62BNMtsxlXjwXpI4
ESHOEfsikP4rmCM0u/08xE3IloI6qT42oQhM4EsFT6T5Lt9VUfmqu/zZ8lei8bHuiRVPbgOBe/1/
l3H6bwQNdOd+4tIGLXuvoHEZkN/8vnnBbGUWeR8SobwYcOs1M3ziftZK4pdCE9Cls98fKbsq+kpm
oH8IEscAOjKZPtDT3oLc8BFQp91/mGn7RaR2lj5u1iRPkNxXT4MfDZHjmWQcBWBuBBDaOvH5maGo
bC3sZQKksnW4urw3zU/4sZJE/OLs1uDdKk+oYP8rXMMWlKD+cecr2HffHNI++JPa3WANAgxwovQO
K0FG6f/ytt7ot7t4A0j+R8RoKTayigxz1srhl7Q+lx5CBabOGxQq4vIAXhrhJWXJd+dvH/KKiyPM
gWDEatpRmC45PRSjMaPfUTVXz9OeW/nJNwlJrtGlt0OR2FUUTFOY/di0miWkH5SdAGaO0lEaW9FX
Ntf7D60neVwNxzxq9cgHXiisUaQbmUTCHFkU0HL6bhJYEBZubCOhKSWGOR/7TsLNQu49KBOzr4vo
Rw18d2rIiE9mCVVbafNoAlTMOWqOmniVjh+WeZVDIJlPWA80vu/Z9TBdQ6054dtsEL75xW36ibwl
Y4B7sxnfUo1UHNRMTN0iL/PSYwpxnwY63Yor1n+0TOLseYF84VCn4F5wI+AuyjKp3Ts+9i3Yahzk
4GE9AY1N6qGD+Q0sClP5cNwkfOazlfwM/Whq2P1/HJMnQhHS+LGjbzLE/elg7mu9cmAiis3YPQcs
6idHfW2eA8jlwa6DtX2Ehdwx57/+gW9I/wrgn5DJP01w49Er4K4bhtYOlkpU5OifBLF7+R82Wi0r
sfRTUUuMDYfhLBbPyYaAoG4Od/gGvOP+6TOnZZbExEhWAspmHrwMSGKPxgD8FkpcKdS0ONB0lEMX
FxrLnQkBPUOhT7ETujlPAAs5R7JHVPn3RNFEbSVwZqxwTP1E7zzRBvynh+DVCfVNHZD8hLR/0gKZ
RciUK2MmM8jrWMXJ0AMHecisBAW4iHz/WxL6D/DsOzElyqvwAEN4Y3Pe8rW1kKU4e41vzpe61lc5
moZ3r198KDsA1+vGL9FO2J1G5jbv0WJqUqNUij5mb7TpoO3ylsJW613hNFc9bMmiZ13zYTiVsAPj
kQZL+BgmIo/ToiGafLnAkN4jrwvVzPCNwp24KNl5SvEcsA+mijleYAe1CtLHaxIVsH1IVs0HsMax
MqRMSdLjxBPLK+9YYTm6VkoJ66g/Q+2Jzd2RlmJEk2XYYOCif3Jd/PPouvKcSlvJhABT/UjyUKpR
PY21CkoF06a/h5XFJl8rKXxD0as+nTJJBNKK0DxaMZ2YdC2NYgABN5E5Dri40vmLGcwkoSQLDDT9
r6wba821L7yj1mzUypGaPjo5DAd0nCTEJXlpTo0JDrkYaVRz8wo/k8JETANLtI48Zf7b8N7kVx/y
loSPdt1aJN7H+rpLbYOzrCAZyA8u7o+fMZQRwT7eipZR9OvMO20XBvStht6jijXEmcfxWqOj6WpM
0YTPmFSk/GVAbvt+RPT6TimQREd4j/J2y5Ks9dnyJOro32Bq+mO5l66+zVQvpX5jSVTJhyUbl1nW
AVeay8U1My3iT3Yf1oxaVPNN5o/hUIcFZQtZe5/9X6N3CGYRr0cZLJT6M40RkaNT6F59EgL0/jif
scnaylzYf+HcMBeTI3GcXhncU8NEC9FHwJVKu4ctsN9yPhuo6AbVmhUXvGq+oc3PROq1TGFEQ/Hx
YgRNSuGJIbS3kbjl5QwGnLG+jJu/bA594g2aL09yUTaiNbPpSFUDESjly2h+EdCNTgFI5f1tl09F
J/hYNRnXpA2hgdyNk5HjnB2m52LYYneV1JBcqt5RSG/pNGxkjqO9YvXqYCkLqWea5E5vIBX59bd7
WQqku4D7/Um985rWqCxoHmx6ORPacGa5G7SI+QhsUH8hC62Kfbjhnoydjq0XLuu3SZRlewWZ1gU7
WE4XrNLHlIvXgV3bSF/lmrUwBrLyJFNeWm6WWkcH+qqeh0CyyvqERuNUWiavBMiYYoQlZSlN5KFu
+J/jA5SX2UhzonryIkDAvREwSO/+CpIfH3/OMJqUb4+IXbt+/JOFPxd9kGUhfe1MIZ57ZyI/M/ph
rNx+DlsvdmLYdeHZqG1P4MwdGcWqci8cgtjYK+1FLxd26ZxapJexm9hA371sogprE7A0bjMtqE/q
2LaksuLtVoPEFoHHbnpcGv9KoiYRqYamXlWL64JZPdY+TLaDLA7tQVxsdJsAurVzDNNmRceix7Ud
Q562hRgiW+wQgVqVPrLDZb3grHybQsDIm0bKHznaikKCTXqoVxrr6up0YapQD84OwCx2/HT+ng8I
rrvDti2KTvr+CARJ1dR966jtXr4/3xFaimYxK76w44A0dsTquo/L88ccp3w+EB1TE4o4gfPSe2hD
l+yQOFhxg1gxNuKtadkaXp61WOi+hVVFjCvttQbFk/5AuQBun9StOygLpC/A381xku2Vi2lmi+bp
/XNDOb9Wxa5qPUCee5yPjTUpaJX5iJfazVTN6ObfQHdi5/iH0SOj9J9r4Xcstc1d83y3YFJXyVwt
9dMog3V6kndzPKt+o8gRs3oChXeuvFfX6FAgrm9Sj9SV6Q3NYNo9R0VG8TeBy2ccMlG67qIzKXcb
E+lx4D9j0Gwewdroc5piYQOV+vBL4DnCUcbdbDv1fMrhViKfAB+3RoDtFsSEixCmZlbAHJ+8nics
YikhmJ5mHBfdxDfAQt7VToVglVZ2qI6/ga7JtFMJ1GAqpUUXrdmy7IR7JLP8jXTEnXmRVMVTM/KQ
UcZTZZaBVvyxrBtwHjDMHYQsHoQU2ccKw+FZsfHKgp/yu3Bkdnq4qtvfgL7bKs70TbUOFiLLS+tj
0TEC2snu8XTYByP9+LSUK+EAfm1ti82sKJRxU2ffe+FIghvo5jR0Cfv/JqxununMoBS/bMUrK8TF
DRFdsB4xw+Z8a0kvzB4UM25bNPEw3toMLwrMu8WoBNHFwvjY5XW3IE/3uEzAj2Fnf+wEeA0xT3QJ
0fuojp3J8rYCHj0rxEo/gGKAVS4apser1VYh3rkq5hRPNc2c01TRVxaI4FtfiFEbm3yuJ+xVR457
4sT0xFX9nOmF/Tf3awqMIcpYDJooRSfBc1+sbSRVxBwkVtucFUgtpZckRlt75gOrG+QRxZcpyrSs
p0P2x06oQRzf+L79+tnx5gYvFhdxPSq8qE9I1g8wyUNHAT6JdlfZ+JSM1wwILIzhwqthRS5iJc88
TjgR07Hr6ZrywRbloHLxLvwG7CAyZiJFB78Ww3btTtbZfwwjL4o8gS3sPy0amPDIxeb36yMq45s4
3qFQOHvjiSHOgp460gCEjN22TuzvZJYfVd1/TfE9/1je6X130R7aEAXAT9q1UVf2Zb12+PsBrjQ5
JKibajntEtTg1ERkb2HA3iQfTYwaahv7AtQ8G7Et/kJboyAPQiri7GMnE8WEETMJPmEvYonR44Rt
lr4OORe/IrYF+MhtnIa7SKbMerWhJecGgi0RvraXNMELL8bjEvfCsjqQKjdHQKG+93bK0QqGw3v1
SP3sHuMXHOcmwDKbB07paJQlQSFi3fvIfKwEJXQsNQpQl0isirfFuFBOocRqIMnr9RF7Yo8xFQkX
lfSP921SS4olzE1zRqyZ0N2tat+gXI2rIKLXfMItZEBk+4oLY2QCF1Im5t8cF5M9HBzHqUV0uXPi
RMMsnIJK/Yt0WQ5LkOi/FJ8uuFLnJNVlonAujcli5GEXa9gxkS5fsIudl9ikM/cSouRlm2cDEfgJ
4rRpLIad9iMlEdGkk3+ow7yDUfjB3YRS4A7b4r0s6fa2SC37hfqU+Ei5OWuLrv/FnmNFnPf429wP
ObsZFc9bU7diqlG502UFYGZHWrWezn6Wxq3YUC++Lr6YgZH3RZbmOtaxU/5O9RCJNzCN0TmLEd6I
js2+ifCLH08TLS7lxzX6QqoKx6yxKPw7V1accdFxL6+quovCW/h1jwsWgbzlZLnm66MWFoFqxkKq
JAcoIg0Jyx4WVAbN+4BP4c+qJz3eOOn/DZv+hOAwmnTGGOmFrKRtjo4ynCesixVZxn5HHCKGy5+N
oo+8KDXXNCY6GHCPch5mc7Uwhn5jqQBF4dRPtUoivHEvHNYmk8co+BbQ8UWrMySKM8Wpy+gS8xqY
p1tOd+oFir4inWy1ZJNl8CFnRj7rGFy7zWA4/nhm2PVJtAfDEE+AEkrA8JNRcj5WbRUU9qRunzTA
vyusmdccn54xQ79oXzfKCk50ydPG9MQxEE/ivh7f4l70I3rw3xNGutKeK3b0Qn7+yej0FVHeUwya
M1DCpaA76HiAH/jMj6I54QcYmsBTf0VyhZVb9FUqINazcUaSVzdCoTNtVz8lmwgmJb1OpRBakkL/
u7TvxizqGbyt6S327x4g+jocKcgTrBAb5erkf/XYm+MIrXeP09zxY1p9j26ziyEGNB6I5hE8E0L/
aJauMJZY2YnfW5KlrlEKAEyeI+q8YcgBhE9pCDXBJCYaDs9EleU3rVOeoucgzV/C1igixvsQE6Ng
wVJw1XrtRqCeLwIX6IzNCfXcm5cqdyTgid3nhRVjoCzMBWpntdfWMUT8Q8Tiwh+RLZnp4V+Edh/A
C7kTjn24olfBCnczk0S8N02eX7zRuhxZe688BbBa879iwDRrEWjDI2slhs+u63MhZ/0/4njK45Qx
Pck6S+Vrv7cSdVm4mByLdGuDqUcBo1q2hxh+6ZBVI2bVDx0vt1wVVmI5W1IgIhm/YSOYlRpFEDTc
b67U5jM/Ks4oLBi13qf8VTuYcOJaimPKL/CjlD+vhuvUTrXqBZhJ0kqpoHAU0pCfUnMS93qIvu2W
/sIliqC26Pf3hge70mU6ye3YAIqtDCdco1PAaL4hD9Sp+qQdSodatGxlgTIY1Xx5sp7Oj0sdKRL+
xdmAZfwo3+/YTeZkwDzzr2UvsaFOz6DwJqdeUVMs91USTB6gVUr06Kz6hdQKSGu5RB8YZ47q3Ign
9QXToysxjppVuP51zzWoU+kwsulj3qgBpYXMcqT/Z0/LOwVf/9fEZWg2qqVzw4DSaCcRxgm3EIof
v/azqhTo0qw56mBUJGQub0jERTk+k5Vcg/yrWwO7j+aaLOVbwG9ktTDhd1wSvmicTPmj4CK1B4yz
tVkdDpitCsXPZAMbyefk6Cw9xR/4g86iSf/VYQ9rgIsHKZDIYzkTzAqxP0LoOPO/RZKZY15MQC/U
h33YBK62dtDO5vYA9h3KGzCkqjfnkaxwZnwm/mxYNiHLoqBqBGG+sAV+NJIVVTIq8Dk3mC8sCbsG
brx7AU52L6DE/YWxt4FpgVnWVk0uSh6yQT5zQZoD54ffxdygV6NEYQlDLAyfL6zyVEkKyU5a/SBT
otJAhnXZ11oaI+GorRr57vxN4gl9G5cOJt3j96Sm6jqG/6fc97EBdLr7Z382x+RfGNhA5ZrWDhNK
7s1ggYZa06uy9n/RkEQPyp1S1uIqbvcT4URX3MGtwti27XW99cU1Yv0q6cW5YZRPbsEvFbGpviYk
QBaJrG7Ld9IJTXtTEUEIL00lrBfV3nMooJsz1Mk9t6CctSeeTFfsJ8t9G5AC5XNPxHMIz5BO5iCe
ULf+ICPxALWtSdH1ZKtqYmp6+P2oWHDVjdyka7Ex7nYGhjNUKzr9k14f6Z4XWiR+BR5Yr8+B0fNy
rJiHa4LMQ85CL0jvJf/GwswfYtF+2c5/Pe5KriwVTAzgQe8vdzLxzzZUYAZl2xc1RtfSgLD82pSd
rzE+txMuHoZMmpzJaZJt95UA9QxJzP6d4nzbUnmVKPXFce1Ip4hoVXqjuPTnmW32fOZdGBpo1FLh
RR3WO62iHZ6ZRUtnUAZ5zdv/lMh8A+RG/JNVZPmUN2YxxjxHFiHdtflJe8Zf01ijqtJFR/W7V7K7
Ttx+sr1gdEFZqduNNbMORxw3Ga64A1oJmcMIfnzlsWgJl6wiMw5TY0JlmnQxdyaYuSJmGfulM9MM
qWUg3vUXrYGtBu5ZzYdvKDb1ZQJSOOlGXZ6lEJEPr2V+IDP3UxlojXnMO5AiVD+vgG/6+p0Vut6t
uUYNN+LvIP1td4M++cLwMFn9GATflaJBSBhFes3tnKb8JGDcLCNTAqtr5V9LglxgbzA+NsdeB+dB
VGf/KWFttGELehghOWynm1qNitJl6qagamZcKJ/KAgwcJa3VTWcDOEXW9nvsdLTXln14n2+OTsyk
Pyyu9WJaszD2P4ufZbN4afJpMWtgKraFv+iT7AB9VEq1hghmHb5oEosY/dCLMrxEfLkD/5Ffn2f/
lE7t8Fb03/7rX4qb3n2PMX2AREwuaV9tmg6cahzVQsaG16RNVOC/63BCqcXmbqw/V3kYLp3RMcma
QSxxqD0fNJbWt3yrEA/fXrkAZHEs4RKJYi4u5ojmCD/P6rjJ9T2OBvQFUMq/zRNnoOd2sVhlry9b
+SiOIWanjcfVcTPnJjHcyy07254kQqnioO6osObMtgpg6p350xgBg4faOZgfoI2xg+0Rj0EexAOr
ezjVNBVW3yhaIH3bs9TEIW2zQo3DnHQCXWf2l+duSaODAyLaWp1nEXfwIFCRgnY+0uzrrClJZ5XR
DeY0GTTfwPBXXSmSxIilPr5EFnayNGjUxpWLCjI28pPZMSBPmPHe/+jiztuNLV0ubw+3s7i5GxBg
Cp0M+Q6Q50cZPK2Pj/QFBpwulzJ4wtLb97o4HahqbwXQRdXKHhBEEwA4nhr4sXHBvFrewIkZ7kjc
hjbOqPyHRcDIUClUOHmAbhXZcdsXBVE0hoQ3r9lsDAju1jRI75fxDC2HWSFXubopwuNaugV5cWOd
6VAhTWX4cs1nlwMU81WytQimk6cEDbH754xwmZmJbUluyUEcW4Yqp2f3MJxjt9n+ulqrtgZ6Qos8
+iHUzxOFz2BWeqH2YTWcpIFj7VoGUg4NJzoyOMs6qCHDTchM0a63DAmuDjNeV6VFOsc77OjM42hx
FomFpVuGa+PKERf/SvAPvsTfR5Sa4jlBahvTKjanc7cRifRh6vDk57r5jy/0CsLwoZN0JC9haSXj
UzrCegRvZYsoN5uOnw+4WEdzz4vTlyhNiNe5RUzLCFa/hPgIXnHKam+HA8GY0hyFxrnfM6c3AGxG
lZOm6DokvFmAmN0oSAeoesfhBysTPQjlNCwQggUc/uPvWjxRcsN5x92abEJoGaCpyvLzbee/yat0
KS6LWg3rVejtIYeLWLHvJsRJqvK0kVN9t1a0fvFlyJ/aJ7JI8YYqct3tx9D5DxUOmVM/+VAY5MD4
rj2MLEI82yaF8sqhRFiFmCa37IDfNSGgoTV2eHFiU0dThKB/ybCyk5uGaAqTd3g+epwBO80t8FkK
99pl5nxqdJZP1YUtgRncyWdimeO0eUNJi1Ybv/N2URZxhKEWG29LANH1w7GsO2I5RhpRMsVitV09
KuFIUmAI1ld+JSGhacxZw6nUE6S+3+Ph/wthsRp6Ukb+29CbuYqt+a9UUvWMVdaUa+RN3EW6LBcZ
ivUJ4GRz25i1MxLag00eh0mAZSKu/NYCG5TOTvcRz9hqKh0fq67Rrj8XlYk0QeNqBgpgSkxge3co
ek85RZ/pysS1ZQb4O7pVWdE+m6ipU1DkOUGS24GYQwDWVK4Dw0oEjEi8WIT6K62erVATReYLPVUz
nmscCaOc8D/yO1gQoe20heA49D50tDW1F8Ly+Zv+FYCTI6YmLXxijzpI//8ib3jqXVs6bnvQra0w
g8HEAopVfTO1uIUKsJ7Cj5asLrVBPM2qXKZAnIcJK6lOKvQBvgbJKefXtwEmzwh00g8CNDAEjUuF
UFJ2PDfLWh0F6h0CJd8EuVrIzFwW4o64OeM9B6XwuLnBk4rY8acm+TVVQgoHnrrc+SIIylSwcWTo
mpqOpVXsj20yg94ZbA7ab7ex+SOaOK+LiwIMNYaq36ooPJuj1YiRNsmYJNkzyCFmleb321L6xlCo
gkBtYnkWIhQthRKRmZpN/JTlzoPPxDq1eTS+kELhAzpiZuY3UB0YVT3m36uqE7otKSNUhm1TNKZs
vW1fCGmt/UAbZE+8477noaG9kZBYZEkByjc/zPAcsXbc+ypMl1lUR89yB5BUIXfoJdOj1UJ5CrYi
OImOQl2d0CUHsSVQJqebMxwb9U4Gzywonx571y77x3yeWVEhvuFA6AE4EChi9Sk386ftUAl67ecx
02AaA9DH2j0nfdZOAOWhkL0aHvPJjsvgldkRTS7aqwCJBstYiRMk/zEEXLbaBB2UOnShNPpe1rhz
UVwnikyYjoFda39JKnrXC0bJPahD/94weN6yrUCmZxJHyXJ4HAiEbKA4wGWTpH2PTgCwBCGnDfRl
Oilc39WzkEiL2ejqzOSHej6rHglipA7cSx49N08ZifMeaRtqEqYYwNPVA2WQpa6pYWc0v0ztiuRE
6Aw4PS9+/7G/VoaAl7lL8QdGe80rFwYUXOqhphwrMZZc1R/X6ELb72j52ImhGnbqo+zkFz+p7G7u
Bk8P9ujmzydOU0WzQTR2bDeKihSUzJ+bLZnWrp+Kn8kqb37M/EVZRAIBKpy7
`pragma protect end_protected

// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
x1OsIDebis699YiEhL9zvVaR4y0ERDNZFfrm/UpG87Lz3GASi6GZHERuml/rG3SmPNo2SbFUvzmt
IZi5K/rjTohUui+jl40jzZNc/CNweraC4gazVlF/haUenF12CvmFqjAS32Wc2L/JqNNjaxiHaoS8
yypnoE8kWIBBNhzaE9WQ9HtaprJsuWhhja0HgGwAqlImK9nI2q8zx8QjNE2Flh1CdTiB/lnzGer3
KIN82M8S2Xi57z8rp0rPFy2pRUcuv1otbIWj4QgTKHGjfn6W7mA3K/qLq/M61jNRKpml6qF1sXAt
Udfn0Yo4X5iM9b2J0+RNp8SlewLwZp3/pRuFjQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 26128)
oF2yha6OcJ5vP98rgOqKAtURxHDHqZhAX6AHkjUnF2RBTqyrHhFJKrF0P22hugkmGsQ/Bvd5Y68v
jfcejCrNcLJ2u1cOTsGHjMsZE0MoWjnTuheOYA/o84roGyRAFPWc2ZtvJnNlomRJICbL/71hjL8t
sPe1ayI8RSTv0xZw9l/bzg2iCKVcbk9gJpRmYHaWCB8KyLcXx5BTi9V9a7zo0r4GomO2Ok17fT1H
cu+bIKV+R/7ndrIv9nJcdulT9FCEGS368dZ/2D6rE2RwVBKquRA1M4nCWPbdCdYGqmJOff/yLfhN
nR8J3fS+8U1AnTt/l3TT7ytd7IVjbeKub8CY6+PEXSw8hjfHmXd69ThmHxMP1bDzZeMFo8/BHE/j
+LyY79yE9NQQeuZJAP6pK73dFS9useRh3ldEFJGXuW2txRlKJfuTQZP6ZL/ZrEXz1vBLj+zNrh+i
7AeysYyShzG8mgraMZ4yQVvijhmqnqtfcFQNux9t9/8Gd3ABN9eWYnveZdyfqP6Dnq7xfZoCMK8v
zhub5j8d0ffylv6T47ul/osqTKTLrhIKKoXJpA4kxvGwVnPfMgZ69Zyg7ok5p74gaTOYIwqcz+D4
sCnycXoZIv2TGoeg1gBxva4bjo/pKiSFBA2oBEFJZghKwD+wMYdTdPh79kkyqe7cK9RIpjrdMAVy
jKWGbk/lhxAe0DEIHJ7KMtYaQJ4KadjWmAChZbRkTBcju4H1+kAssCIOIKgXobcoKFsx3aQgN7k0
k/lkq5iOYhycbbqFtCYEwRgQtJTgleD9oVSeRvbwvjilU1DsYB+Fdq22ufXJwoL75XoF8a3Ro3fR
a+GN5fy2gd5TzZvwB4aXbXL1Ah0nWxDRYWUxS8zuGBQtmTO5m53xYlYXwjF5hwOuUCNXAqanS+6V
r+LzsGqFSQNVpMZWHN1fQxdpaWgup4AjD2z8Fr0IxmgTd47l4LgXnnUNsp49/rPbM7JUfPXeP5U6
osYmRvFpRIR4wDghgMlzTVge3eTL2QdSyb+UjjnX6fi9BU9eYciklzAQyUzuv2vIUtczHhITWstZ
hfFRkqymVCEVAaAQnfhEx6vAeVuukioelYPE1N5EkGulmOSkDQpexdxdJfwrLJPK2FXYhQx2kPe/
sfcS6HGZh+mrCF6t3eZGlRMEr5MEX6rVpc7p8iwlTx5B9Q71l2rtt2porHI01gO308LVown04Br7
EJSxDteyssOxKHQwdQOtU/3OAberiDt7kSo/e1YrCDahATYMtNaLl35VMkyX5kKfaFhkSN2Y+mqI
9cawx6FmZNfl9fUho5g8iQw4BI+DHSbN6PKPGZIOi7lCnQN3P1qv3Z5vYuJq4lw/Y086ULneLZT7
CIWPqp6c0+AZEGlMo4I5GfD9KwLcUvHtCcHzBSkIlcBXM9pTPA7E8VZIIrPJ+PHIZzqrR11n+dH7
eCfHTtpBhvKiAjZgBjls8KX9mo67DegRrFfTVK+j0s0vaCRF3PYvNMgD0uywcfpWieZTIRUPlgGd
YcDmgdOZA+MdXABYvhvxneYbRLz5Jrtv3bkfKZCPXXQDCBAwCtZb17aI6oQ7utEj1wraLT7sIbFR
P9P/OtmWPHfku4v3i9blE9NggUdwcmjgLg9TXyv0/+0e53W3/qQKJDPOHdQLxBs9n4Ak+luKksZo
jp9zMZ2AmodhAaO9tmqbNM5ZQKdIi50Rwhq/T5OS19v1k3Lov9W9hhkFO9eh+RaziQKgM832fIcn
Q+DGxd3A1EZ2SXQcA/DSEbHV7ekUN8RfqLRp31jmlzJtIpb+1RbSxzaMzdsm1MXQawZAIVtyc2z0
hpo6MDgUocAvSHJePp5gs6CgxKR69h8g2y1qKqnzOfWm/WP0k4Z0XxfhyIOg4juHBwHDzUJqd1G4
Wyths+IZa83opKWWm4Tb0ovss7IR0pLp3zGTvdWkKNwgRElR4OFalae2YD6/0G8KFkSwr0Be2Bhr
VMFtOSbFzZrxPPb8YoeBHHNnkJSHqQ5Qdp3Mou4k84hcjyPZm99R+1B58jxR30WQQ3tjymGJkUeO
3hKtPGUpCQTNCJnyFSh0/yzugzdrzNXAzCasmjofDmuKqJmxkw9iH2TkNZNgHUDKaNa4kFNp2CZP
VFSFOElk6B0e6XO68rMUpzwBYFHwgU6f5LNiyvltjDiQTCMKCN3S49ZcDIRUO36xZzJaZMIK3qW4
pRbWBynw79VbTQfUe4ZYGe9f/qVkQXcjisznYwLtZEZsN4MbJgndrdxap/o5F9s9xT8N92JyzBeP
HGckLzIYOhQo9Fjl8SDEA33jbIswIxig9i9J3GgecoHjv3fGymgjSkBM2BXKC1lbQZHmgH+hwcMo
uT1Jo5AZDG5U+TszUyX1FZw/TnS/kH5p7EUM7OouFEwEm38vRIIWM7aACwN2w3NTNePZ/5pSHtR6
+DDeS+osqmDWzj614pr0fic654Sguaybcbsr8kVIWgJLAMbTbanV0JYJ+mBQaJZNp5WY3u462p2I
oehpuzXQ1i+xVAzw4UHWVk1/XI44Anaopc0UvAXUmV8kziYAE8UXhtmY4unEleVY+rXgtb0XllTD
w3kOKs+r0Ubbvm2T5GpzZDGtSr48MnbCbsUbAMuocByCPnzcy96ZUMODN7zw0qO5rHf4RhOSnikL
YRjj0f1TBwLCJmLd6N/E7cBCu60x5GIWKhviU92h+rx1FhTpxwA6ABoyNwkZc8uC4+3I+6/1Uy/X
NGQwW9R/5NNYe1aLiPEbbNogGGLkyXZWFWZka+IXnSXhsCagC2pWrRphA3cdlH0Gh6nLOsSEaQXG
oveXZ9KZFz1ONaOseBF9/9kbHRXwnp15spdb2eG0bdDHF7PHB2+kx1imXYSWQkql3D9pWJ66uSBM
CCYsNW3kef4Kdw7cQR3z8aYGwhQdCQBwRRIxQyFl3g7BdcHDW98/I+mdfD+4Q51YkgnaYX6ncPw7
tSO9tECExvCFIsDmCeGEJDrTEaYqQ5LS5RlBPoelGdY43GnAn8T16kkX9vZ+nOL6M6CRtmCroHUz
0/07GtA9dbGnDWYaDxwoA1IefLynEyq0l6Q3FWUr8i/uERKRs9liMujxyeI7WGpKksg5ABQP4X62
BrnSz6bX3Wtzk4Ba9BjMKG1ydGEVYkn27WY70RK+btBOmJz/4tSr40ZqWqvEKBAFAanB36NPYXdJ
RomtsdK3Qwf6HOSOiLwpbbt+rIL4FEnNxjhHvkBDwSwU2spP10n+zL8I020wzp1uDIYceZ7pNkiG
S1k31U8OFrQmhDJVAZjUUuIJuGhXOAttbl9SrQdv6oOfK4FU9qqyAKRWAmJtiGvsU4TQXQIlOoQp
aVdhXovBPNBMEcjWchEsshTslCANKpOYFlvRPrM3zJYr7vjqgBhQRS+cOnEjEYWrVHhi9j14JZmO
eKoltRtY2UCa1mZmIyDwrrjv0aEMlfSbOIB7RNLJ8l7RLZ6XrD9SZcLIbFACwGna61L/wDG/MCK0
kPV+79/Zy0pfvYCwcCQ7Gc/SypfPywLrDzbuwA9a43swMW5tf77aeJvgGjI6ORh2ch5e63wN6Rae
OsY7M4x20XpgiDwh5LiDAj6pqMn+Ofxinkqtjr8jddBuCg0ZhThFExKTuH16vMd0+2Vvn5CSJOUe
lx9kcvCdqQWrVg2Fv2A3o88tpCOWZcs09DOq0ZYGIZWhA5b/xMznTl4jEPMHTlb09K3FXia1n1m0
50yPI3hEgSN463sp2odm7hkp8V0Rm5q2AoDKOp890o0b1tHpbBOW/1pQweCpNEr72xWeMbstsKvD
rE7mOp/+Ifbu4kXHrBhz5YgZlq8yhqMDm8l7Lx5sB0V41N4mbLDXcCfBvXAStG+JUmvI7jfrkViC
kS8KnpJbWznXMa317wtInymZG205A+EF3yPqDDz1qbmdPXE3SRZ9VN0vQ/MLBok9Fp7Bc08LSSVJ
7EMwUgrmY810+BF7LYeYuNiC+YztGJ8UODTJvsZVR062KBkXDl0V7qwv3n+Yg4RT9TvuO52xMd0z
d4K2v90UN+/JJnYopGPNAT2W4mihdQAcjWTIgolSoJslQ5H805l4JxhW8S1CUJ5x4+RxYoIoOjC6
8hTm4jl9ILwL/d7fRHTUwFAEFGOVrSEcS4sTNwvQtPdlm70nrM3bVdG1g/8cGSar5EimtyqU0jQA
/cReKuxf3n2iLPCInrw1TLT7/kCcuRLwB/n0HluxuUhVMSFMSn/HMCbFqKuGvdncaTrMw9vWH150
U7WWaeDB2VtlYu/qt813HwJteClAh54n1r//FUwzzzA3CDpNbptv/gkhJSKf0lDCkFlKBD9IPrx+
GOrVSOPnWUTGFJqHy10E1EjAo37MXHkPZc0AhbJzgiwUyJ2NKlTKQZ4RD5mwJZUumKE2trhAJwVN
zIyzYaFcVN9P0CiyFSuUo9rPt2QgZ+Bl74stKXUtH9TzmHEwD94E1b1Nr6AhqSzBb8Vnz7c6zR1Z
JuSPemL3Gj1r/FdEZfYA5T6kArAXKmImMbMbW/UvEBnMpYz029Snq7nurNjNylWUGLUuooEvHIfi
muNsUHZMUxqabKPyxWWtInaVExxhm/PQTPJliGRf2OxIsX46il0PsO2dVENx6lpK7prXGf0vDGO5
yqpo0csLwAIXr0yL0a3WzYTUZXY4Fb/jmc2GCpQHrcUxEPl5sVOw4YYWXIykdarIBdUVkYFrcLin
tV6+SHna2DAsZzTRjPQIGM28FmvRGZ76kVg2vZTKZqn7rK2VZw8R582Y7dZeQdOUlsBqjVcFgM0j
AOOwxkLtZXAs2yu3w05nyV2vkTweZW2AukcyQS7XRKc/HXcnXDLQpHeUOF9PR3cq0Dtd41fTvKu2
tr+m4tcQiO9UODk5UVU47aNxUwIt7nYVNhp+0WYpPPzxWjU3s19Wzc2V5dSqgkKhuxgDq4n1T1dy
FgyRJngx1XOCRI/YzjMsRQp7pcriT/wGP1EXV5Jsy3s+MQ0bpJoi3PK83HU1Kp6gfJa3Xo02SCNA
LnAcUKb0rLjjue/wkTLvQF9p1rp903SPc7Vdeg9MKrEKTzz0d8xPemq57ZFKvmLoJD/vGlAU/YKW
ACLXO5SMitserc0+L0mQz2IYfxwvQPJaBCVUowOr5WmblXtiDsYMs0QeD0b3h42KU08AsMuPgK9p
RasAxgaem18xtHx69pobjWsAsEGp7OsyUZ1aOu7ILlH6heSBBoBBhxbp3txh0qipiTr+HJXH1Tqp
KPuAvcQ+euXvi0f5pPKrCwW4WDLVzzCZPtxA/zIGBUJPhYDMzPjgCTYgd0oU0Tv83f580Agw18so
DSon7VjYmQs9u2hfv/KoxnG7In9Trv1+PnCHTKI6tldDv6mQ0zSGx2HTMEcqSgXdKHUu1oZSfeSF
wvPhOEMueY4UsTymRxxebqA/LMWfKQml6j9YxVWDZtVH8GfWgnVMufJS2T9PIMW8VwFoKqMStsXU
W7DVypw/DC7AQmRMal+j+XoX/eFcOSxQmQLL6QoNjdWbxQ97n12FKiUaS0F0DNEARqa8tiQNxCpH
aSpRrW9TLmY+FgcA5K57/vbUUoX3eq9uukf5obDofP1FyY72pj856esNkTuH7ovqm0FqsPTcJq/u
DxKK4YODSW1zVR9vB41a4rK894SCqKNuYOVx3bSaW7G7YNVooexR+jwSwoZCkB8IoNwFW6SSTdrq
YMOnv8KtoNIPNCBqDqzlz9v7dnQv7V+jRzOkEA+BzkOiehq0Em2SR7h8BU88skay8++gfdQX7LE3
SmTQIvnXT6zLtpTMGDkFZwF23td7KPA1Trx1NixQcZnYONGAR6TOvLki/8mX/nND3MoLWCq2EAUO
9SLPT6/M7gWbgVq2WrGpcy+njwiO6G6tqwZhK/7am4+5/aPxCkFgY1jmlXUkP/1gz+HFKSbpEz21
6tQqlpEFsdjA5wn3hTMfemjUeG/NyrWsjVm1Twb/LTciaeagEkDz95pdJUUB74a4WKPhdTgWI2Zv
8+Hn+gDi/L5z1bmd0ZNtiJ6Fv0/euN4ZLlyHcfNQdqNNtgJhgkTS/Pd/aFyFz/mOc8iS5cGJ8K/W
6OEiF7c/qVQquBTsiWWblxgSwh9DgYf2PkXyae29ja5Ww/OBfr/oZ3t+c3pdmlhXjfrYtyYnYDkW
t5+aeXQvTA1fIHmRZffoflJ75QfgnRXBMuXxQZHuwVonRB+vnjIOnf9fUHnLdgNukY6Dees8pwXM
ZegVNUaSblnoEhNUUUXqrQhW9/HzRCHq6Tm+zhBzbJGez7Ys7RfkvdS/7fyuM7YWJYyPqWMsfyyL
9c2YLxrwERY6MV8tYkdVrFleTXw1z43xqdU3Y2r5bwYxbt/wkYCi7CwHqKKCno1/birF7As9bLmd
rRG+Mh79iGTCuTNus05rxHQ1zvHfBvqBT6n+BXL+NVEQSG7Cv0FTxSDVVzAfXT6Of7lay/JO4IVu
+Yw+rg/WsxzpnV0aR+DLiMKrDqipniqr1uZmKcd+eqGXR5viR4cDhkuVxRq+kyhdGjwQ2o2E+nqO
6qW8JI3rKkjgnmTosr/E3CneY8SsAQOZbzzKnFtXAoU30A2PUglbVfnIWRL56rUUUWWWZTWYssMh
LHxh1fsvtiNyi9jFbftudOa47pSMdfYoVvGQIs1wo7l+ZC9q8Mu6lJ4ymlGrR9/fhr1dVoyqvBgl
qVr7Z8Kp/7d7pRaKaSHaWMQd6d6xu+usB5/INhAJQdApGpcdUQ97S9uccspdYuroyoxUQgKPZe03
OWXts8wS6tRCYdTNLi368FwAVMsHw1I6kz4ysM0KnGrIhZFub61/PMBfp9fdCnxqtHU6/h9+c6l+
aSnoybCh2+8qXReCbsijo6T6cOeTQS0G3JyYo2MH2QnhUpJxoMT1XHMN41ioXjuLh1dArSY37FIN
43ngcevVF7g7+wPw3seE/OoBC3cosuCNJ4qPW8t4Vp0VUeEhftJH/hfJTr46Qgu7uJWUQOH4s+6s
zAO1Fx16aMVXSFN14dFlfzG4sXESBJYhSQsdZhptJA+Z34bTEMS5nSMgxvuEXLp7vQtlZ0t0huaG
bWJDP3LGdGKsb275F9JJhOS8GkxwGXtF9LY+YCEhkldC7XTZodwFNeSIl6hG7qRkfngGYvK33376
JL6e2SrNhj8Xfktg2eK4z9t4XPVisWA9Ys8R3ys0nu8heR2fSkISlrSeTI7Wl7NpW8k1oxpia9lt
YxtZhC69qJtN0Zt5EEaDgMChw3myUr1vBdujNEvhh3q7prezh0WHgEHjHuEPTgjZa5hep6Bfq5oN
pJIzYrq8FWZlahjozJ2D1Tqb/5owFAfgPHaz8BfYsx93+fFLms08kL0f2k83jSe93f1ioxjKdvqk
sEHklUP8c+ur2DnfQ99EZb82N+FTfemwKqVAdFXzXoPQoKqVZ3OicbpHhMCSJAvsdWfsZpdA+2jV
SxAIls8ykHiB0H/JZez/NQaA8zo89gYgbuopL6z6j30qsjYvtffJSTAPo/7Wj3s6A+OVHeGjLbUz
3oqdLZWsElFZLzCtd68R5QfSzgxt5t7ppUVCoNai7KwZahsdNQ0E7us59ljPEAeF2IxhNMga0uA1
PtaAopVBpLj4eEXxT+x29Sc43x3j3F4mTinbWgjEhzooI17s5+2XoyLBNqn+So4bdLPKAhdjvima
I84BQAPQ2HxzhpuzZndzpBTINvfprieGsQ+hW6egkFSTIAT1M9Hbj7u/rhS1Tq6Dy27+FmHxXiOi
aIsTt4SxnokpDPfYopxeWfXa3dIR4gql3ZPFV+vMHGW+QcoQNqVEcdI3DBuUmqzFy/3CJqNEWMYX
T93Ivt8/tRaEZLRcxFhKH5dXITQpKZ3m8SOmNxt8Pl/V9rWXMzNXa2IXM27mKiEV+07SEukGbQnS
TU/I9hXadR2BUcB1NX7T1dlQNAUmO4Tba1Js+O5lHpjIsN5l82P4rBks5D87ChUGuGzTrTRYhF7/
gHizqrVKhJK8/8r+SsLZ1Ynyy+DIGObBDhy5uTvpiCtzR06SWNbKK7gx6e2xruFoNiWd0Clyciih
U4Qr/4lmNAd2gOz65wpN42bQ+0yGqRP0JoIDnDL7zEJbcn8Efm5SbRlLTrWtnJ6JWV8fsokSGL2P
xe7P7FVROAqZYJCnPYRzwEPf0dl3wRxqHgCz2DDvgNcjkuFPo+hM7xmVbi5e5ptS6FStaAMsc4g1
CFXWse6onk893Kc75AogANXb6CiBqDjvN0k6Wm4oQA9xYSIg8MWupflIEkiWUxVXVKMqp2tXQljg
w0Bu0OKQvN1HECBIXUOvrzeTVMCe/NthLB9FsSG4pxamKVIAkjRFj4V3SJFE3mmvNw9Qd+XP08AX
4RdUtN4sE+dNiBt48eK/eD0PXgNDWpIjjZal9eAdugx0dtFqYSOxGcOzVFX55CVQKEE4X9AfziLN
kbv08n+7BGArmYqqxPhIZ/orTwFRG6XwsiMsB/KDf2CXLaXexSO5MSaZxEgTiACLTgPznm6ocPwo
EDIguJAIqUWa73cP5hX5qTKis7rYjMK1VPKga/YAg6pUlxMPLJ8bNJc7iuaEw5PVOBuhhwTqCTKA
fJ6Wee6Ir8MY8AP6XdX7TzNLZVBjJmQ1SB0WCUa5gF5FyHPIK6pWUL8VnA+1zpQDmpICTnTyvU4h
fFdtkbnu8wUz7h+0DzE+6SbzRF5pPS9t+DW9chxdOG3lCZYEyRLQeNSYQiBLqXSjgIZtpZB+oxZr
PsEWZtU1H7mamKVMJFth1813evHfiFSe1n076CrXUNoPM6gzOTCEKQTdaw9sK6EhZrFaMxntMsA8
h+8cqX3QQoKHIMCF4z4U00hNrtJMk8+V0dMM56GroWyqyqTSjyms11hpHlZpj0OXVRTFvw7mxlKG
hB8+4d76Vx2MDEk48f1G90Z+6FFYhPPMtL+MXTgcYdVJdi9/uYbZZZNPA1NkejUN5HBrtlghlHC4
j1JSlwzwH+ZPx63gsIVAf72MtSdu+y33BFKoJ78eaoUM+D0n056tgk0qCS7JqK0SJyw5MOHmuyEf
0pUR2lrcq5bOMHeQjAFF34E7dM8J8+FXWblS294/5qeCmHGekdDoQzZU/S6Eh2NBQtl2TYE5o5oP
5ySXodfTj8gL4IZ2kL/8lkUMdDXCIk+ZvJnkCLrrSHp7kRbOCMjkeBdQIHtgSVoimaJXk8Fr4HgQ
ZeYZ5HHhkry4vAzYRn53GKAx9LLGd0YUA/8Re1lfrqdOBdDHezoyu1gNrm7UDECyVtBTidjXHzmr
i9lPpxgwIIUxlRqokdkshH3V2xF1jlA2Q/AawGRxaYbWhtfGdnD9NwrXlDrKBWMjJhlcle/tCZj/
ebM4/TuWGGac4BdFfaNwO2SqHGRM5M5e9+hKqq1Zoj2BLEYCpqGf0k0DTl6cxNrGsKz+Hr57yEuz
XTJBjzr+BpenAb8xADJf5sGewfvyT9VqjfDTSjtSUTqQZQyoCkbWCXzmc5wuvicnYYV6dVumtVnN
7PWUoPl8+U/GSOuCqQp0eCk8uqCcwFE7v1FWqfPnD4VPotoPAwEYC7ZYGiCqV1A+rFyPtRaXnOsd
/tBc5z5D5QgNNqawYfp6d5PAwDri+obEz6CU1MDidnPqGV0o/ThOeZNGmvZ3tAuAuCRYL/Jq3TnI
KIbYMq/sMrtJeauEqA+NnWYLzq9iAftlconrh548neGZj6YP11bOAgjxK7cMw0dupd4Cw3PSN+Lf
7YMYXXn08ML7lTimX7UxqCLqQrEF0K+W+397aqSTGDC/u0mGKVAFrfdyESdleidUUjpCtCZM1jiH
1N3r58minFxQgoAudNLzKj+mz7DAgsGvSOnLNPT6RVuS1xa5x+5nvZAzlzWJYWRzAZBz3x6geLcw
LlLsNzL/LGiYY40+pCP2PNAMxNTeCtRlxAhfGafwr/eOVTvDXQNdxKqYRTrwwjlFr1Pl3NqzfL0g
dBEZ0u/IDMiQHSp3Nm3fCyZCAZmo67cBaeWgKNydh9drjktaPzU+vrW8lfbGEtnQWqk+8dagq2gY
HGkmVDfbhcBgZ7zpQUCKDX58yu2vExxhJ+9gT+pyMFlhlSWlZ8bMP+YJtciZ+MKWlOQ6e+Oa1ZiI
0F7A9kN7RQefvv2X4XORlE4TVeDuKbnvrWLFf87IaHzLwQ7KMD5gYR64yePcZE0LsfAtF7QKq+Co
hZrqpZOZkFeXWNUVPo37OtJO06zMTxEZOhbxZcKvAOK81osAuCSMejuOepK6i1Sz+1y9ilL8ZDF+
YcFHDa/YAtsTMyHXC02OvjpOzmUD8ZfXr2JatGhI8rb/mLfytHWsyQrnBfZIOIsiYjIcieygzVCk
sKy9EX3k6VZ69SbPgHMPN/pu768nteBWUOJsgqETgd2dfsOc4y9aQ89B802AJUBwNWN4UGy2qUzI
LVghECz6hWsSRUkTGnbPyz+z1/gotJ3ZsJAVif/ddjNCvTXoKzWKiZ9//pyTJ1YhoPYOZAnQK3Ba
bmPAhBDG1JKMB1nER4EQ1HmDi3BEaPnFvFvdwyl77DK6MAiuykdlmqaOZ6oZuvRr/RcXtTaHwYQI
VifPtR5t9U8bweBpt2bY/CWVPq93FCtbeOX0t7da4dhuFQjQI/oQ/PkF+IDCmecWozqhQSgG9Hhd
DhSLuOB4DU1jjMuiNN8Pg1PppQd9ygYbtiUfiLx/bLZYf2T1HCNYqI0jfNLwNfhouGFZwj2Ajgvc
BE/Ut1TbcTDUfDjXZX7BXRc9HQZ1O4lPHDCienM7eYpDOTxTzLqYRUtDWnm0Ew8dp810kCAdvza7
vxChxAi4zorkSwrTAiaGjbeZZns5LrEKaUSulI/T0dsnYGWzuJGo3Xs5NMRi6k0UwAaopTH/qNBe
1AE7sVuFmIF4Lb3QWefBz1FDKFnN07mqoFlmlFt2imOqAtpZcV6YYwnl4R9OnRPzLoa2k37euhdS
2D8lx6CqyjpJgdT2tT+bq2BGFg3Lh33cy8IW3JWh3g8X+/JszpVC7u57RVbsroP4jimzu2YLYR+n
Eu3sbXirAI6bwQYzYHgNQ7oD3WcgHTpJnyXdlqMw4kf4+szhjWzf0e/aB4xehob8VYVfgiuLR+3V
YuZAHL61eJiF68bp7MN+zbESfx5waVGtuMWXRWyICTh7gsIaAPUBoo3Fv+ehcdFt3Jbxd5Ko5Hzv
A0+3+bLBwwMqY62b2seCS3NH0nTYLFGPQFgICGw2gg75OT9h/h+y1ivvk0b9JkH/y5pCnXdN0ziS
Bhm1kfwpKXGlJ23hqvB0Od2mPm6fZh+grV2H9CwgXWikNRGpnSLH0U/Z6BcBrZji4zCj0ETKDvOG
qqJEdxbs+ibYC50Z3qQo+oh5+PsCKpPmyNccNAr1mJVr1h3adqs/tqj2p/Z49bMep+n45KxRQX78
NarGZt8lg7f1wf5fGxCDPhlRoGj3pwzHxEJYwHh0CsiWguPMPSNA7+2Kdba4hKQBGZHJrNQoI8lP
1Crl1zwY8p2xefAYq0cG0T1G5wtT7YLL9qhFNIJ1y3Q1yr9nzEyfOFMEpXRkHeV95QV98X3EvLLr
XoQJdOauvKZ7VJFv/7xp/swGeWPkxxigPDhBBV2Z49DJNHquGGhZFOhjN0C9tSHTh61Kdhtqd5xL
UeFoSXKapcWLIa+Cwv1k84TJdFWrO3zTjAko9q5If46E168Fo1zhqL+Zrjk9EM48atnr6W0BU60k
+OqMnqYfjeaGpX6L4dE5jw8A8XtJ18S/1C/um6Zh/ZZTgR/SRpneSQEInQGafna40VkJVpNq+K+S
zxm0YAE72BvZqZQweMs0Pc7RKNqDL8FU6gNfNpRI9zj2RJ9aBFmPPBe1hYg4xksmdFDnn+53dYza
6bTj04x2IZ+N5KB9FvdJETdWdIsWWztmOcjxghSODS1MZf8o25XCYx2WLSVHZ1RHEpt56G8fWFdj
J8YkOyt7liWlJzRmCMo5uUtbg7pgCyVjlhgDHISL9Jcc4Yrbe3bm3cdW38YVFp6UT3NJ3KaVetmE
s/haPub1GyTKPmOUZcFnaIY3t63FENCgUSu74FctdrIuppZTq9EC0KoyGqeiik7mPC9APCZPXbzk
KwJcaZH82NcsirWri52avuL+k/F1keuYSga/YJzT000h3Sn8kKvR2UOEe5lwF2gtskhtixR2R6Vc
ho5MVYaIJ62dD90rnP1GriNk0EtG+IQYVX5QPYKfHLfGBPId+oFQD6ktilRA7TAidSoMktHYSzqN
auiQunE1wiXqlCgalrZh9WdaMSiQDs35nV+pFc4OEupNd78JlY0QxexWqlSQCEyjuVOKeLoRQjM8
UxieXGz3DGlVy7xenzIHo5MEEi8G3M+IhXhP+uUCaj/L2mJMtSZiUrm6It++pLHpGAyaTVAFU5J0
RbcSXe5ofN+ZhRg95asAWT2Texk2FQ7LIYHTH852zeKuPTDh0fwJBsDETXs2uQz96GlGmPjgGlGY
s+9tNZAapGnwebOyZ38pA54yhE7APASFxaCYXA25fKVZdXyYmuzSVv6j3T4DRAgoMxEpr4waRoIt
4ZEFg91sH1Tb0sjx/J2S0bNnwGJqWfnaU6ihuu/auhztt3u25yEz84G8dkOg8Q6tE6BiYG/EwjW6
a+Y/znkE3s4PwumApro+pXWhDqvpzvY0rDmGusn3BzAP71kvtpRaC9GAlO6bM6Gsoa9G/ftcC44N
x3Nv8IkoUCZzR1XvGoyIB5XAnzhlRTdgjuu3ePVL6HWjO9P5jeYWFvg1QVafZBYpdObd44sxG1Qa
dhFidRGW7F3WODLaZFCkFyPrgP7IA3qp0kf70Au+Q2nhGq19YJpE3rTiVDvbq8gooNV5qTmvU7j/
luS03O+GrYH7F/FasVHFbbowArEiYp8ptEf31h6guIXIeFkbeUHL2Ew9VSLTfwTGag1R5ps/APbt
5mlKNMPUGhmeWY3jtTKf1FsOtKE23932zSrwt7bgUjV4kV9Dm9Tiiraoun3QsUJXz6F+0nxjZwLH
+uPRa8W0q5Rt5KPoqhv3Alv002Nn/k3eyaNTM5jFT2UwyETepg2bb2uOYLtjWfXbMHTO3TAE5DJV
gNaA9Z9s6O5bw6i4wHUvv1AcomHsPzdZW8a4ZexfibPWmsftjGl4iMis7/3JCjDdm2YU1SZhAkEP
MeX8Q1TVX1lp5Tr0dgXyy4iSAg0Iv1i1ZwbYWRDudfLY/MvgWt+c5L/qhLDrU7mpC9RpVMfej5NL
8qTgLeHIM+1rn4nRXqBjj6/SuzhHVrnGHStT2Age9relyjv0eYoYSF4zBGf2BOu8s9EfaPRcvd9A
NyZKAB4F8pn0wl7aJT6nk7sAX/Z9GypSlJV1mFXfzjqAq1lY7L8PI8teL7hnlb7lN6PWgDp1Ypci
tz5nPsNLdVevFTtqxY3rp3VVg44tgndyJCquIgMgeWyeV7w+B2GB6IzpZKcojSJqyVewIUBczjtv
OEKpNPf0N2HLgVXeGXXIe4h2W9tLxi9GYeBwEoTcV7U8ZjYMgxYMbPfqrZcHtclYnIKAIAwlRVvJ
+KpER3NqZivnb7lkNYSUNn5dmFDA1WYmMCuemvky44f5Rk2tNgoaJI0p8ZkK5iXdl8MuJemSF19X
4QgP+ycgLhPruu9OmdwhXIZcJajG47ke/EigqQtY5Nbg0rfobVWpGvOcQq2lWz8AcoJ+5hg7kVxk
LWryK0WqWn9TmpPBzB+xkjACLaBma+Kki8VXfZzzUsY4+LAsf19wczAGC6fJP9GW9yVDvzIVqk+f
qmlU3sc2A/hxtAhPGMO9VDavBMHAzhyb9hcc5AGQnlFYn/uoJWXjQFRB2tX8UmGV4FKZluosgKy0
+RtZ4VZFilT2VJsbXZEJ7Qe4eM6td2LBNjqKLp0+BwqdbdErysr1EjsqlhS3nFzezoQecrKo/lYx
4GUSVGtXrK3jGPfKkaYofQCW5B1lyW73jxc/I2ZWQbdo7Cll8wdjY7vY4sZiSuC7KL90il5zXpmb
HqfNoHJh/bB26WDIx6vdQUB/VqasFO1DfV7CYCWqmlxHOQ3725RRfD2V2xF+gTpi+Bjzd0mFrWtk
1SsqMV1vQnRUpsTjQIWFqPclGAToCAsOoHfjuP3UW6J4HH4sumZfI081LDzx3NyJ1ZjaL8+TsARk
mcHwEDiDJE/17vcsL0B+y9DqeVw5tIDCJLwVEbbpcQVrdcSSfya2rmD276D0430jZNuhtDcLXuDg
OKQ1K7nk2+4EZT6/jX2vF6Zrt0E8699v4yMqJWTKg6bZagd2kuPTkN21aYPdvec2nPKTtfznHRE5
jBySsPbg4Zbx5DyX7cbsV+j8OLC4fB2ofI3qv/jCmJb7D8twVHfJYfMb8CmKn6eL2ZwfI5LGLheK
dtQYkEvVpOf2Xlkmz6TC1f+CdUjihogVEtjPiZiAcpHOo78mi2MAjES2tabs+gbYkIBkhcirInYE
3PzA8rzNkcfP+5uqBCqBHj00iRhKHpnKz6Jd/1Y58YLgfrhjUtWtqEXdnCDd5yGm8oA+zkdEFUTs
yKH5SpDFnDe2JCZF6JMmR2JobbQ5XHv6CZPHzIg11QnmyxfJoHt53rOP0Kcq1ilqQIbWbOW5Bfgy
zUKpgHDywwpckPGDCo87xwfe6y+GTO69nDdp17ZElXhjDY6qZuttw/SQ7aKsWXO49zkorfKqE4Uo
vjli1JWxjDnKSHyqVhiV4DypoIPmadSZmuKiOAJd0h5XJAXbv8oLwahIGjOX+3SEunBGz56+VcCS
Vzcx7CraX5+9rbGfRncHD1MBIqNLeJEePTfTf11QuNfrqmCO7FclbfotMsGlrh0x7LvOgyyiq2il
4pn4iLtYo+kPdqEUgb7CVcpowDzHepClipLB4EfoZmAuXaSI6S7CbpLmQinhdc3i2MsC6pNeuPYE
0wsGNzfESlvNvmR7WvN4BevQOkHDX1yYRnjqh7vN3ldRuaFmKonpnIkXK6MSil6CbkGTIa6JN71G
w03zrIQ+oG0M0ojSjfclz4RRn6s0Mk//U2nnmTp629U7O/1GNP08Jm7vC0xl+DE/uCYF9eaTmpUU
k1NCDgLef22ihR8LM/tNrOdcNxm/zc774fo2lxlmSvyRswdB/vHCAc30mlpLjjpmMNbScHJ8PsgN
FO8/ltQq0no0l9Intw4j1AoT6HYX1OsU4BaZS/ImW1D206Vc6gzkmPoHQS0Q9yqj5bUJrAHBupYN
sNThuBrbXMG+SUlU66ZYmPA2k4Mg3tWwIh7QWMoRfiGSdtfIoB8XHX7vPPPrA+xZcuvhcO1l7nXy
+lnmNgU+WXYhu4e5O+YQdgULn5CvsMrkRxmcjRm3OrZoKM6yDE6pM52t+Wnzib+QWeBCWCtXzqz7
dL+Gi5lnlHYvj8O/S/ZVtYYfwqdk6XidEUFHobX054QbaKZbPzqrPqrLXBpe/9ir1KaucFAFXRKH
vXH2+FINsP3yaPjvsBr1ZBB3PHjGF10LoZ8sv8OE/SAGALBT/To4GslvHLlgrHRRHmnQl2FBAp3f
9UNCaHYLFdte82ShBW84N2aeJXgztotyIKqBoauyOEWheVR+hpL9HIU0GUZwCmOGlSGou4UMwj72
3RlWUx6lnJThnrncj5mKSG7QgCv35BOl1oKB+RBynMx8gPCjpizo7qJc9A3j/bkofeQvW9bFqJOJ
YcJFktpzTN9ePaClH9WphZIyLc99d+afkL7fWf++7y2Z6vFqnqdMeZI4kghpr+3Ywdl9yZayjVjc
5a57UhEgsdKbqgqophpTrIDXmLQa5qJzHWI781CONMdwpuIj5D6al77wJj9XoOcE4ZxbZMXEaO9A
scoodc2MhAbYLlMwmQQZsr7KjaV8h54ktEVI8sbTkReVMmaJo6UXCwBLSFMTU2cuz/ACMWi8jiP9
B22jlj9CoIu5P1nKXSuAfrKYp6JwKHH+7ozOS3shJ2aeJ+aHVCuOifMzFwD5qyhdnfnVHMQA+JY0
BnNvWL9GddS/a6Y1HBjjz/R+zXy060AgiPKcBxIhAvilk4ZRKhTOf8X1IMs4/UC+HO0FGhLV0Bne
m8a1gqTGCRJz24AztFuQFY4cIRMmYraZBoeGujf36tjjAATD+ulKKMIQnw6VxUkXcZk5kn8dmLhx
wGdZle6gum9JSrbV7wvwCsczgGhcSMUt6beLQ2fQbGQaMOyJZ+dl8NidiGP3hWomEYQ4cA3kq2Kr
+DBSCIpKB/ScQBrfRgfHgrYmClFAWpKXTbWaJXYDtxGwgYYqFbqXzgbr0tRUq7upyPWMLmXVWS4L
+TE0dCiyXLyveVOZd5CuberxAMksEE6wv8B8EmBBLPKyX34S4s4aS1CkNshVjv4s9yf2h9TaEBph
7D0cx3KhP/FTG+g7TFkfIyw2JSFDEq247We/r2NALlnDqstfiwE4YMAWT3k6CcCHDKKH+5eptpUX
0SLSM10tocuwbRjfCuywaaXQQ2FJRIKqXj8G6QJy+iUmKasgv52sEonuVLJazE270JZEECJIRNAC
0L82cipgX2EgE2aj0opcY0X6xwR5AgZ6kMd8igPNg68yOt3kWQ9adMtPN9HlPRKkaZjV8v5Oe9lI
xKGJffKtVs0oKNdcYybGs56m/gGDSr6gkhI6slzkupkE1J0ls8ywepyZ2cNQTyc068uyOrdtfo7/
+kBkpPn/g0nCOLuMOXpOHQni6T0WPKLySRXeNiYKepPXX2oqP++mydd3+tYwVecXw5x7U3lJz3CM
LICsvZ/QOK7RwygxLR2ijPzXHfBTz0z45HZ8wqgaP+C+mj00ZAojtnGy4br1nQDNwBKbUG1Hs+mv
/5sU89Ev+VWRjvtI11mGxEvjv3OX+u4JikAp99mChiRk6Y6sfMq9fCbp55On85sDfhdyVytKO0CI
ulPY93+SF5gM4vTrLRfqLRx7EPHzn59h+VUIfUfIXfyPVK9Df2eG47bR1A6drarz1yPNl7d9FEFd
ndDsXG8vm0XDV0X/mog1VX3JJ8CXoHkO69GgO/9CNTa2X7rdHqw1hLN0fJwnkuiOKw1hV3tw/6RA
0DJYOPqOO46S1kM5AsDzdiQMvJNn8AzdnsoXyoEH5GMoQUqD97wBsrL+BwGiRnSG1tq3JzvYf+Z9
1fGEr+PReg4eQT/VU+OcEloccxtTtCO/J5CXBHDIpuz9Hr5Q0RyLqqSp2zlOyFFCcVAY6yathHjr
4+5MWamAsvjJMSF5FQ7uQ22sjJBPZYphzH6+BfH6wPHjdqRcH+O4HRdPtbJcPCYjp1LBcE5j9g1F
+2zxBFCqM41ePDs/kn9Uyz1EPx0ukUoJfg/Bpn7LvmlZGNocokik2fGp0O0nmT1p17EJH3DLTklG
L4kfRl+2L5sYM4J6LQVmNEnBrs+zK0vri77D6gMD7uGOCSqwyizwqW1/Gb7EdnmDniHMRPcw+dXp
0sJ71rYN1D37DPqE6GzuL2cYKhOIEg2wwaJhaU3qGhoODXQXFGOWIsKIcUceXfLrU4CUob5oCIPA
lueECol09s4e8NGBSEl4J5jXS9UmgXUJhfHoVje9mBZWXjpcUZPBCftrckmuQOdWue/tqzMQWyP0
PbpE3VnAb7JZlWJqZPelcg7fF/POVX7/L6HU1t0Qt/J8pTbNRkHjm6XWiv3NBmNbWjJNC1qj5n8W
l+BgIiy2bVINMB6DBtiDkbvE0Z64IK7R0UfGF7nJ3NaafY84y1bXkN6WMmckCSRtUtXKa6MrqYe9
4BJH07PFfbY/3XHQbsTevfZyKBUVsnJkSWsIFj6UUjAaH6Cnhm5zkrh1URBPva/oJA8wSWLvbt+P
H7YXXBZu3iYsMn+DI4ZrmlfTYRiF8Gop5Q+2UUVLjUGYla9aJIGgSzqwoiEK5HZG7pW7/f+kDKHv
30vhcsdG++J+Igl+DhhBR2ZrGfzxssc0hNFaBL9gnKdYVSF5oCOFeXnwyN0qWLIx88tUU3TGTNPV
tkcOT9yPFnXvsXD0wnpyg3JDGOPl/7E9bSHyYGgjT+yMthnLafbtW2KZKe48wrYZFhI1ECwsvYGV
Xxkl2+B4Njk5NBHw5BRznirINOS1eK0osi/s5Q+JHMRgb9o+teF0ls1aSeXmyeuCNyCxc+C/ZT5R
9+xsSNFwFchRM9wlz6BAMvqsfjSBo0pZ0K1atTSj1wqTJ+gTVpXNmDh1bK/ps4l2u488zGje5t2i
5sdbcYFqAmHMYbBlkv+/Gdk7iDG9c21ct7f0B5LzU4u931jB5i0ysyme23ydo/i4KbpKy0xrEQP5
FSFum0fsYw+cI59i438bZDIFKez539zvWIVMrFC4qzLbJcRKyYQTijcZZl2LW9H1OT9gLNMXl+9/
Pr8dagGJRqf7UinE7XrIboLCkMVOrUfhCj2TpngkZ3qgYv+3QanaTWpvu6J/YFuqHzT3ZmQ8zbxz
vu6f8mrpmnkp9kIGdKd3ZWMXaO29ssJSh7kyJ+UqsGUAMqiziKgwdwyIz7E0VLMKv+D6pqDez7w5
THU6BLHwVVW557OaLvtZDX0HbjpSWocgRsBxEqiSn13HOec07YjEkFQ3vxG9wPt7tWLTLvrI2OgC
YgaqDZfPu2gIAv0fr4OrllQhvPiP4GkBtRpaPGaZJMW9u+9uzgUMc0hxq9cpv7LN9J2uAgPd4XNE
d1g3R1c1ndoutLmOK6uJs2NjdCeFo3GmdXYSt646/Jh6OelVzOaYhmqf/JCHNmClK5809SjJMzFZ
E75W3OKtKJhLkSaJvNvipK2P0CpSX9O/Xt6Ij7QRznCfJZGLubUTPs6/+veRknUi3Ijw8E+aCkUp
6N0rDa2htqF0DrRaMdkyYDcMZOZ6RsIbvlmxhAvIRjtFccnGA8X94s1hz0K+aqRVaOh0jAZ/hQu9
WkNQ6HqivCmgiNsPeuAIrAr4HqQXISR+ClS9B7sO0Hgs9EsKGzMNe3nEk0ZVVny5gJv8EYUqjngD
AcpO7yXm34iFhkZQgrNxO6YXruBbihGd9xSu18PHqtjjLT1ah4Cwop8RK9lYvIcuH4U07tMfVFj2
UfxmjEDdg5iiTdn/+hlcBKGGoewWQHQS1rVqFoqAd+W/zOmxlqWZgvdijBJB5Os+UYMsZTLvP0SZ
Pce/9/jMHlrnNLyNzoxwef6EcDrpFQPs0nLGAi23gGYkFYQoYLNHDfwOfF2GALx2Mvajt4gLT8MA
5evifD7siFqOhQftW1dGERiYKoJwAQ/Tf5meMj8Db740onfgvuCx+RNBaHQAdFniap9D6DdhGQyZ
5Lrd6XRS9RCuHY2YrPSw8eXL92HqJL86izEZGqOyT2wZ1s6HIeTrUBoisOV5KxqvvKu7UrX5dGDt
4sbB58xTmqlms1weUsAvHMkRG/3ecoYBvRTWe1u3AR+DDgh1JNrNLUbvhD4D0S2Oj0nVX6CJW8NT
f96exEU7i/qXOT3wp5MlnLACnQtQyxWmcAg+uQz19bt2fsO+Dro1LtqMdqOhPWe9o1TuX54IVpgZ
c4WXosX7HoevJQwwVktWt4kD3HApQseXzvM3RnDoNCZAKI72Xm9vFe3BbOZOtbdDaF9o9wVTjKKh
uWDGiEgYaO37SAVg2r6GH3XMU8bJNyg3UcVEXDQGtjex97kcwP/I4qKOWVEyfRIDncQyNTKk1Nff
lw9h9Oj78kUl0sA9DZ8+SU6yiB0JsruEGb4P1jJ9TU2OaFno1EZiNQwTNIwzePb7JDrTMLtOvakT
68Vw5C6AnI08bh39EJYlOJhSmhUP6V6HhaTmRm2DHH9JlD/mj3ZbVGBLhs6KxGr7sSfmQminR0So
9ZfOOLrSybbSin+4Ha0c+Y/FiblqdDgIVeVnGLogW8ASPgZUV0+tZA17uH/hP2jdIIuj1B8ARfin
ZFLg877s6CqBQncw2UmRvMneIgKjbFv52ZbBkDlAWl+79n1tyIknbOQ0vogxVj8H8JEiHrELckcf
tKzIvjDMrjwpmyuakYCRlrk0sj1PsgMg6QOS5cRLaOWCKWYmBVk+1DsigUmTsh3XIurhSY893I8M
0uRSArQBM3VrnrkBtRN3UMinMueguBalHUYy5sisXhC/MyA4bkJUd5dPEj/2hmsUfjbN/pkLsK5t
DLseBBKhPmX7eLDmJ/ptH3G60Sad96AKo59DhKdmAie02Zd1tl4bk968X2KOKqGTCt26nurWziiE
TKd0TgJVQ681gXinxn7n8tvWc0imB2mkQcDMAIfnLCsreD49SwD721PqbmpD0TunNwm4sHO1RoVw
53MLOqjh92QeuQJwoKOGvPeOUFQLYFIUqNGAJ+NTW8IyzBJAx5oBwJHaA4H0ZUb8vmgbycrL2/ev
t4oLm/hLCUUZp7Yx0jkNUSA4O1qe4YhgvZFDIbLPfcB8VtDdHhOXJB24yLMfnGPtIGvCCJwVKiv8
SDHFwwi+GQkWRCM7R87zvdNny2w+ziqVH/BJSTvTe2KS1xPQLzoDId6lMQMg3qMd2nQxAp1JYq4M
cBJlxpmLj/1c8T6Fl5vHASe+5hq6zBu+yxx8UIPO+AIGzuOVoSTkbebz6GXBGVmGViN+N/t2Shx1
26VRucvDye82BIQRxGisSX64h6GHlkrocTR5M/eIaHqL0xUeuPkaDePnHh66nmU44vXUTBs4tVum
yTPR0kwnSKOTEE3rkGp4yVKOeUOshmGldZaxPLgXwPP+lIbXmt6LuaLaHDKy3GlEOSKs7vJIFDMr
05e5/wLMxHP3XnxN0qFN4NQ1oB/rusWlvtNLwwPx7jEUMGq+w21mW5+7CE+rT1Iws4SyGxIHk8Dx
YMuylWJXcQirUdFK53B2T06O0OI+twlNOCqWeo8b0s903JozKRzLFPjmimKkUuWbecFgnAv8ycuJ
ohCea1WDGK4iBCUQjPyK9UpMS1hLRg9+7+A3Z9wc0krX8w1LpIiTghg0Atk8fYx7E9/QZIPWdtPU
4w14Ri6CFE55cYZQkT0C+qcJMCmggW+KMQAFAFZiy9Oao4bSt6tNkWj4By0xPj+1fijLjeA9+enJ
SyI4fc2dZbKI5DY/dB1pAGSNlLLLyA10GMoqfWPSJZjQaJnEBv3f9J0xCgitqS4/D47an3mcrg/a
wxEDLjhn09GTidEuzlztSsgS2J4UYJWGJD/Ex5Sp5/lXO+cPg8Mxj5s/P8/kG3PTw/8sJgQbuBLQ
S1dtYqBO1iouzlT2uymydwC/w5n4jzsVUQP39NnyG4VR9/oxsTqy/nlqZKvGq4CxBgFflFto75IU
yzb2FSZX8xfIUzd0iJRslkj+P564oegk8h0lKDBGwfN5GHAFWOFNkDRpULTOZlDlXqvN0vZU3IvI
xq5LywZBlvNVaH0E5HGnB2N8ISJs2XGGkg1kZ+9DcUXHTpp/ppdvcGek7ZF37dVr5BXe2XYzHWh7
5QfqdPi3NGLMOfjU380/tBPct9MQ/eApnTIE8ksUgk7QR8k03VwPn1+M4gM3a7W9WhAWdslL3beE
EInfXNa4xji2I7FoZxrp2QTODbkNMgBqfOfS64bS65F3pOnw66hZJBh2FBWAxpTsj6r6/DqnxdE/
LjBJz2wp9dFy3MC+TkUctnr1cgTIL5y9xpQYBsxXPlcdP9DRw8I2Bph3nZ3nzdOuvfbXrjA62kxI
nFCvSTxHSpz8IEtQCQSb5PM6QON1q9b/bNqVrnTxKxoR69lsbF8fTTMLKAaqRzOmoeKiYVtlk359
uLgO/srEYFKEBpzIh29S+8CZmGWULHpiKUug0s9IbRgwSvbH26E8Hsxd1BxNKDO0PCSU8Fnp7Qsr
lS7Lzrrd61SqkygbgDczRyV83sYpg3gCv981p0Bl/w657u6JsMn/cUuudnb9MkNusGh/R9xo1T3r
FOz8UBjsjXmneEdewAbyVyweotacA4LJ4+o+hlqTvOQCGezqRk9qtMrK3ydou/ocFlmbV68e/D9y
XmriLgb7gTuiqwLMnElwypSLF/IVhwVl2HKU2w06NvZEdLbnha43xfdXmfCeMl/RGylfnIe5wXKE
uggCnlK6/pWBTgiaBn33SgbfAgZ5MTSBSgDz0ykr3z7ZpVxAci1HToLJ21mw6UOOrwWyOs6hbypy
coZXzloje2GlQnVb4JbCpUifp5Pi3HQnx2wwR6QiXXkiwjijVxeL7PJciuAA96jHgm34pZXNYG4p
TEQ0ubTR3YEBs59GEm0uwf96qK/z8W0CS3nuPjcCKuwSD93w8lAt3JkXH1lm+loR7CB40HnTroyz
GZaxtlXmIVyGtP+96dczyECw7WepU9b7gCjNKtSNVon85uVXfcZkTJTr8RTt2k4lWWBKwzzwM6M9
WcQe4K4LHYQQXxG9I7VTwVQf4Iwy0e/faM9W04ew4aRyjzBcamxRLopy48lsxuIymB+w2IdyNQoC
RprWKZfX97/rV2pG/QVaQnhNldRoMZiJX6VOkRhmFGnrYV8pg5UrfJWPa5QopU/2ItveX7RSQ9f/
Mee+k1Jv/JLz0/0k/h/IwpBzXGZ6FfrXxpXzUDwxVGhwjJ+gmCk/YzuGo52Bi5BUOI4jxnj5Veb7
oEZvueyzd94CFVT1HKMoc4FHl8KRxwNSX0JDMbP1OruxNPRulpFtZ7FnqORNqYE14XxEjCq2vMVY
Og7k7mZAGHhAXYQ6PQd+bElAuCxF8Y3veEfoiOTweDCU4EK93X/hIPNLVCldbMpOn0tiYmIJkQp/
LhQUuZqRrgnF3gF5SfiVwW64NgLd6rFCFqXHHpBvJpHpMeYBWhq5cdKwr4aAPVjIrtXeKpEd7fhB
7an2qIkGgSWRbRgwSOVeTmbitj75mgeGS1Vwz7q89EfUdC30H8J/qD86UZvDUYFUIxNGrbbqLhzx
Zlcc8tSR6J4xYRcXo9WcQLN5FrxN1E+S8FZYajYlDCb/vny4zX35dQUo6gCmgJUkcEFhcYx6I4wm
dmbimJtBRGX+8JodSBk5j+hWMawAiSvqqMV7PqGxzi6JtZ4op3ZYfBatEuCfl2wm5F7KaH5sj6Nf
gd0uYcQ8hhE3qN34XNqdCnXtFg1+0FvYra6JKgxV4W0hhyx8RbnaKkZGMOCDDQgm9NQnbaehywUB
VCLtze3NCcQMY0iIzOYejEn2HbEVcT75FzDXi+kgF7aETfB9eSKXdpkxhpH8118td/1AG+i9syaZ
LQdZnqZvuc4i3UmWcLtTKM9soy02GHXqFaPpdC4TbmOMjiVMbgDpmCimkgWqxp7mh60MmThUIA50
rFfYiCjtoVyBrU8IXgcaFv6Hbbyp4+nSwFAtHh7x3PFm03IPa/EtmjF/VuL9NGUrQsJRl53pPC2e
4oSY5psNwedzEPsA4iSIILi6jy3k15oJXIAVeono1n7vYuqU+cFYHpMT03yRRWM2+WFLJzGuSXjQ
XcCx3LFfEJHG5ahqTwpw5Ht70s0jrdP6DeOth4Mv3lnXGyuHZzoFWSOt/ZB8sFUzS+7LE0cvV7Ic
2vudv8XiINzGPx78tBfQSCiFQtkplD+DMzazZXtg5yZLLTuGw5oTNj1xDn7GN9ZhrNwfLHxkPHrG
ZaBdYR8wEthPPOMtyeiXmid6x2SiRjvUf1PQOqzV4sP/xpD8DYrchksoK6YWKWn0VxX+yCHzro8Y
YuYFqMoz5yUy8N1589DP+0tRQfMHXeMOte9utxSmxdYZRrkXpXp3KvflprWJSoKkXc4zc+LoOb9Z
FEhRG5zz/csXkSSsU5a+OXxJOa2Ue0/KMD/VdbQCrH9EUfr+EciqwcEHYOEBtBFUExVNQrLm3cFs
T7pHmly6SDfomoNCoZmr2fwJMKXZFyFSdmvJj3aWvqhnsD+tWrq8RB85KpiZciJ8UUZsBLIfy3uj
BksggZL/QEgk1RIShVC2akDx5UF2sJl0yyZGdnFVJtIYIKdJ7U63Ua9QpOYzTr0x6WS646V4mgX2
F1yK8RP6PQO6aIpq4eGyntsvQXrsN6NggPqOANL1WxmFP5Mxy2mSOstu/YXcsJFU91ihe/bEz4IL
0Iw/HcEG0OSMj63IrvNhvF+1Enmc/+NwTHvVrDBQ1EtuaWpQIDCcTtec1EUYvrPiwNEd+y3iwK0z
7FOAvvdZTaZ9LnfMdoV+8dhhadjOcuHshr9bhSxxnVc+ehqJcBL2kYLzWh3bH/jgbk5CV6gTBrq5
Lc4wkf3sDnaMqa0tR/eC2vyXQxWdF/N6Tsh0CEPCGZWg2zkEFiTyEW+PlnPH1Y3SfpEQzKzV025Q
sqrn0dtkYnQbH2hbbWJtEbSuvH8b7VHZXHq9uZX4kLhzKkkk/oTAS9ncB5rpnxaeT9SS5Sm+7/Zj
pS0KnxvoENFbE2FYlm2aRoHzi3l857HlxJr/JQNS0TK5tzTUqYu8jUIzxRU1C4udYFGqj2uNs1ud
OAxcPLrsEspgyLePb9pQ5Gy+0W8uiEpkpPoGpQDcUKGL6ShvsEWIvpRM1wong+KvIE+gnPIShanR
nFUqD2jdwfWlOCQcRvZ93S5drR0NKamclOQGKoIqco7og77FleXouKlhcH2wj9IAlCOGrhRh6E5S
Lgm3JsUzcmpee2vvablmTBeYwOu7RF/QHkSq2JMscg4IDnKving3s/BYXfGOegFGw0d/tfMGnfzI
eFj/INpp7HoY5IcDa/5rYjkJ26Jfr5qbQw7RSr3lywOcjXglpulWn/UblqJLnwn/U58dn6dleY4h
TCOpuErBOqL+XZO+qIlvzzNU5quY2VerzfBhEkR18AOpQ0oVhTa8Z9CBPDgc2nhAqbHG+HDwTWju
Z57EZDOSl+zV7d6NIbHTeesrKpLjP06l720tPe2KWzXyQS964qEFzy3sra2EdNM28QsfPNxT8Ody
J1I3FXe+6f0umoVgLx+VcXm4H2S0DOiG8nXraH+ndr1LalXG3FBVpwWp3wEzFn0BM1YVPo/9gJZ/
rINuUAliD/VVKVrgrLQCKRddF3cy0edarpGIhOXfOqsXYgn4PQY8HL2K1y4ZtFib0q2Xajqp8TrL
12QtPatNxM3uq9jDLUuGNViEvpDh5CKL+UYL7+zAvxXvzlWLBCSy86PSE51B+2uTw+tvrroA5IpE
eSgF0WjLy/EKwlfvEFm/RaFX55ap0TMPGMG56XB0fX0oocip5TmqdcgrNbktFaTtsbe4NXD66za2
BdLJVnT1QpHEKpj0mvYJe6J6pQSFdcXsoUJdhInOPvhV2nWdc43Q+8xPTHWC1iUl5rbZ+7KEXII4
PSaaOTdDTay58+J8HCqPdMSikN8e+qTkIQrBpRX03nk1Wb80jqtz9I8CCPP7DSPeuuD7RJSa7usR
X0j+IzT4vBJnpNR23isF9wBBEeWh32FESusfY4Igj3UnrS5dGi+crXvt92OXX9fnlm+9+vxLojzN
bO9FTJlKTu9B3Ja7PrYBe3ETENAiFCk5fhjYp0AC3gBCT2crfJSuKTcYZir/cT7ytQr3CHzqanXr
SgJlrojJB31t3UbOYdYI4+v9f+EBVWMXSdE2D6pqIwPss5mWyuJSa+QHLH0kHAVqtF42cfC7qsOV
WpZJ+4ZY69p/U3D9gEuEnRLa2t3buwEIFJ0+WCl/mjfh1J2nlJ/ZeNukJ5wLjEA8nOtkiOXWTDr2
KhDrh8ypM1ytXm6s4c9VD+awVKCB3sHhLJMqWiUrDoB10EIP4SQ1eDCaQwEpLzX8nSLVFNtZSF2s
3nHhrfAKDcehA1tIxlIngsBofMinx4iG1tCOjCuEstE0ZtQZK9I9zJMXsSFOnKxv50a9KhEn9N1y
qwX2hRIjPhpxYO2JU5G/uJQhbJd2Lc7+S14z79Bm1UvIx5Aa0b2TW+4vJY8C+T6s4WV70KXBsN2N
aUsgAqHhv63Z2i+60Gu6cKbw5bE+8MaBAhN6X0YUoQXUW8DjbFcGpIj98R6SAWbSNmVeCj7ii4MS
S6HlniwIHAgXv4uT3sukZqa6VprxUUgR9QdDru7BRllbLCG+AKUtzUzg6KztWvP//C/fAtBDv0ER
j4li1WDQ1CYcu8GOWTbp8tBI3OehKkPyNipwk/Q7C93dbZ6zgVenPKqGL3ldLo1Ac3BIcrCv3p34
Z8uAG3lr3w9YJwkSfuLhPFUVkG83LUV6A+K4z1Ou9dMZQdsGEJ2ko345tOSCNqVC8QhMnKGxhjnM
HSebD+nQY96RjIZTmPvRgBAdUeUEBlxZY0LedHRC3RANqX46pX8rNXfZZ0LcePC6xcqhy5iSmcFr
+mdtCzFtMnBULxZjoBVUyLi1A8uaw5GtE5i8/z4U/k6SbcFbL6FEBxd2iaVTvihj60L/abNAIAjQ
hpzvQG9+IvvmNQwES7EcrCL6teVQ3mGVpW1UMF1J9SUSkaA0cddSdWPaCXWEzjU/P/0WaTD69jXn
X1Mx981ldkmhWPB7JszsJzmUxStlavmwT2QuNAQiklg293N1W7dQqOVY1PsKXwQsUl5I/Gju+IGf
sYZpj8UCQ+XexCVFWYICsok67FeJIpn92bOpwTfRt1A0g89+rolrvXhDGCXB/bJ17Xrl3/6n3/j5
gRgAek17FnfL8FNYt7QKNA4ZHUSW0c4aMG9N6Dd7Hq2WXMrD3xHRGe2Z6Y1w5MLqyqsihnfzNb6q
aABhBnb6l3AIqmQMrd6nznVk26D2Igi6rOYem2elbx7QVLqH7d/oRhUTRMMDy2zlrCPd9JwXhkTy
LpuEyIHyo1HlQWUV3IV8T+ZfnmCKr41tLRSdfhsMf2BxOzoy3Ivi89uaTl8JTjmJHcl+LgjU0SAe
dXKht7cJ3RpPFiHMRuD5JEneagbIuNjWWyP2LPLmdTdJetCVGRfWuN2OTtaPox76hXv0EKTd0CeN
xzE85lY6rKGm4LmFNQ4XPBFH6QmF2DdM/oZoHRs9jtZ7Qy99RhSYEYnPLVCNGUPRaH1Eg3QdBPwf
c0CmxIFI9sGl/Zlt2PbcTPXOz2vdIjhpRcQut76EHFcSCBe6udSlWHOFDI+czU1Dv5N1MvXW+cvp
qipvZeE6LddpxeNbnNhnBPACPEtBRRdpl5ftAZQVS/2o334OJReEdpzRtFSDBlC5t58yhZQgjpLJ
89WekTWaEYyKnHSTTqRfWiuvix182QuE4Uo/P7is0lMcO4DGJkOsy2bifuacWQNF2rFd/V83LkxO
PdDmFNIMSPBGRlIv/cJQ6Ota8A3r2eoQQCUB0jqX90n1OYt27Y+f8LW0opyU6V1luLjAnFUqQJRB
1+ivKf5V/S2qvYSE+AjSXfgbIaKtLT9D1yVYUNqvTNr0iJ+Iyh+sJhCm+/WyYg0PMQ/eQKUZ9Q0v
4ycAWRjC5oOdGNNwWrJbGqO1GfhKv+MR79SFUU2Uq6qRaRKgELdQigc6eKFncGdpTyVRC3LaxZpe
IsLiQhd3U3vLX98uvgrcp1dnKIYGsn7MaP+gMUHc1I505iRmt/nmWjXlDM711CyuJWcF82nNlgQy
7HYsG/BQOLdKbH/l9GdYIZ/Oz1gthTz0Q5l6xOlZqvyH0qzMuZRxeixPp96UfsWre6ecDr59bV88
GlyAH0omrc4LCOZYnEj/y/ZMwiukM3jXf83H6ABgze3qDspmYie1ObG0pfYjC1O89/WXS+2RJfHQ
3L1VDjr/OCKf06fMezq/Ekq+cjO8s8IbqZUcfJ160A8Jir0E2iVryY2J/iaZ3pjdxu9KeQ1aU7Bi
IfEx99q1cspE+YL2MxjkXCLMqiRyI6OH3Dku/3OIu0GPheHgghqQbxwLMAr/b6dfquusrHaAg4zx
U183VKKZu45NFsaUZykEoz/7iStBxdXoh0BErXu34nvFtdh0yeGfmk90utm9bfH+ZJ2y/AFiic9l
CpeWhzYVTGKZhnAY57p42VlqnnbOMEBrQ862kUaaKA/kafqXb2jXFyEAuTA4Eql3k4JJ6mbmCVNO
O6zVdoJWknsscINSloWNPuIqoP/m4F0QYr2bZi6mbgfypNcEwnCPo5aYBkqxhvBUOPyZ+hd8Um2W
Eo+bB6UPD2HAk2ql7CXNhk0MWfv2dzxYxu0Ta9N/wyqE7zPzYBzFv1CuaOoqMEEOrRBm8KxdYq/C
RwecymXv8Y4iznil/EdpbOi83lTexeCXalXKOMaMVPa0u2NHD8CCmvrL64Vet2V1iJbCV3OnzDoq
7cJfrobOr9cBvMQakGQla4nGyH1PRKUdpzg3lVhbdWc6eikWgMIZqUjHlcCU19AN878RMhxIH7UW
OjENU5X7r+whFMWGPi1e6w2HYFp5iraNGmmmIe8MS5LrAvm3cboJnFP4s0NEq0X8BpxB1ILPwJ/R
KvZ/PDX+3wfrD7fG/iPGAzooH7SmwKKvDl7bl37NBEuBPmTzRKs3g9HCU06x0HsZqEDxlIcI1tNA
/Q3yt+9vC3H52FI02fgY6x6gTDNrdYk/y4RaTpO9bkocYunqH8anzzZaK77sJ6pwT/T5Df1Jsoh0
dbe5cxGOQiOdpkdlFdfaUDL64e/ukcjRI/u6l1Vdru5UsUf79sNkqgrQZ6BJj2+wx/FtepVwBuuP
UnUfewppoIr2zELgeeffCsBRPdmuD28xOWov/R8T5Aqc0/CP1TjTPNVY3T/aW+XaB/nD1GF8DQD0
Wris6OPg7LsJ3bNJKJHOOABEA2rsVYBTMlR6o0nohLdu/RbjPTDqD0wlCZR8iNzJRgAx+gJFS285
G1nyDKe+rLjRtdu5eCtsJRpR/7btOWnPAlPvhPJGZZy0Sf/jNKvaQDpzMu1l8uTVy9YOzjpq+zaN
yDMck5c4jYP5sFnjMeSLQ651WLnBKU3UoExEQtrGdC+Gd3A5XDjlX9zqX/mgiGIZzUS3oatVaH/K
Xz3g7Mpneq3SI6mxxapU4khy6dyYbAMdptGUKgxYNqZvS/pOAfN0WR/TLmzDlC9Ra7R7LuE9EBHE
SM9sV/C1Mj8zn7+QFQor+HFr3bNMTTLiIbJB9g2d/sJNAj+s/qlUVUUn+mvVmmD4kJyXWrGeCW5v
j5aE/Fr9PCERimpI2SzeEmUdjXsNDSMo8npijHiBuy6JZPXdtI2QMjjuDHrVQQQ9MaAGPbuJjxlo
DOZowYP0rgF/xDu6MBYcso/jQesDm27zdajLplr/nh0jMDN4lDvCxUfkTVvQ4y0l80moZVVhr/zD
z+Y54cw7ujmUjo039+T2gmd+q8FU3LBwqCNzjTr5qZXKEkLkf3X37cZN3UcZwrBCIcrq+1NrKODJ
EE+zbqqg4d9nlhvo5wX6DQsdTUpMlFsmylnaKHdBh1xS7L14iulARaINiWyg5HJmZb11gdlWP0Xw
WV7Rc0A9rUqa8t/fKV220aQPgqZRrG4W4gjeTf1Mzey19MGtX2PMBKjSOFvjizFPVl0ljGo2vDj9
iOswpx6eg/ytYlO0LiLeIhIKmkDgDQZHRVsoshP1SbIJA9aDoRgOmo3Yht1pJGLPPZbEYq0U848f
FKwctD3QArKP78jzW02Wi5xgXkEF5ge7e4T405R3p0TX+P7IsaIaYLU36x2oZMCF2M8h0sKxBE8X
MHrIKe5LC8gjG5kQ3p8T2mKZJ1ZuzJXOAd6racBIv8mLZBMZjF/06/UdTqx+f++UFJZgXMStx8aX
p2PC5hu7yQmPdoD31MHqYlytUSTsGSn2iSfL4kcw8MmS9GtkyMu3BzERhyS/ZEL1Cdjnf3VdyE+M
DUYJMFZyTsq5bKx4Odylfb9nkBvFj1CFICqUTPi89rhVczhBTEFfEwoiA0cJBcJrvX/PxGE/faO4
Y1MBm4h2e8s1JzVWM3/3do6jZdi1Z9swJ1xveMqDqEE8TsezRZNO+628t+322qwKJ07CspZcBrP+
cLnOCxJkpC2Hl2BcuA4s/iAQzipHJpmGWOABNUNiwil0OXdnqJ8wVt+Cq+O19HTqQtt49IZLxxrT
SOK2PI4CWIKUPJtnUIOdU04MLaEBWGbpq6jICRUDVM05e+u3NIyW6OKURpZdPMEnqtksKNhVlGyn
oiItQ9AYLYuLHyEnf2960rJoZT6BQO3yFPvZfRTEgZbcV0OY3uGu/0XeJgpOHptGdoWg6cMI3o0g
lySMzRMWFxSNdku4a5BJqjJ8tooLgy6De9zz8WBF2OIsqFUJsmgtyT1Z4/cQnJWYJVSk7EDTDZ0n
PgGIlIPNB+fcF68G4jBipBL7qKNelTFl+CBFH5fkc1NAu2yxF7NgkPNogCeAPWaoOT04icABvezB
Wb+Zd6UJSHovsPwC0XYuENGd11rsgOeKUD1inwaUzJuVgf3IdHG0OoqYBld8DIOFpViowSuR4IAD
BFBapYakUVv0xorTQ2Hbb94gL8Gz/iJwpcc1W/w8AgNYc8rglqP2QAENp842NgDxC5129ArZXdKr
siSbdDUI/iW92bhpBAdAh8PP7a8qzJWXtT13b8mAo0zPsiqXGUz33gjd3yFKzytff04x2Kmp7znV
sEsRJIVzMapepNqDhkVjqyNfpcsyEzRvnuIyV7+Zq7mQlH5K/YeFdoekZ3VAIpvOqTUKWssOHvKL
OyGaYMvSxHPHeNN5MYqt4fRnJy/pLdOgfVQ9H0tuV0L47aWZcLrEPdL406wNkryMguJh70IR3viN
owno8arAA3i3ZYM+6kUh68KFzPvJRhQ5+2BtqGkNs2e+K5Tl0iUcVMoo/BHXhmD27fHpiIe/qzBG
KFK1HNIA2TiqjpP7uWui7TZOOnaL+hAJlG1a4azQc+EldqStZOlslSwOEMj/RDg9tTdu8oN07D97
pWp3bpv+pQrQzGRAjUZHQsQg0Kxjn7MqO/YwLjUkP7DwoXT2qM5vTfyqWxVkZrMoZMZMYkR/wZbF
/uwo/dS3ofQGaw8Y7WQbFMIxuLUyQTb8LKgvCimWLEHHR7VyYVVQrIAIRk4d7ULv0lqyT3M5Niq0
lPlfDulQoNmqBQ5H2DDAZzMf3BsIYPEGkhfFWe1uRCKgv5K+38WHsgiqW9MdgoJ82Dd4LtF0zNjF
W+ebgmjCHSOeiIyZ8CFI35e8M7V5W0WkeMNRwlZhfrsVPGZn1wvh42DvkeLVhAhxf8yUpFay/4VI
m6UvP5cSlQOng7KNpg2RMX3PodzjoB1anIHqiWqDQpcwjpIzqdSgN3XM5/YA0xKcWBCf7n47PMPG
AShlidGrOFw+oEebhLpa0nP6059FOzTESgT6vPUwop3Q3yI5hjYlTCo6IjjT/aZDj0UyoflGzsZr
KQ6LKO4VyR1XX6KJeDtOuiRxi0V7y8Ex9kOLiMQwPn+sx05vRMhYRQbKrdwgg0IkI29/FiugNQiF
z99DTMU80IdNy3MvAlzpA5pm9KIbbJsmyubOJJt/IrqqzI9laxTlxg0DiU/dYPucYf8/rF/Oktty
ks3ZgvjkAM0AHdBquEppHJEy9xqmw76Rk9sTXhnTURjPeD3LunplwiaOqK04/VOR0ZKf3lB2bmhj
l5wJdyY96JbbRIivwyvDzm93xmpUw85jrvIlaIkuDbn59KQWv+NUJITnUNEE4iJ1q0d5fZHWUUfB
S9dN7oLBIcFecaYm30WuBy7S9uXYhs5+4x+zV1e2v8RPbhmNoJoTnQvCS3N7VWEU5eEnGMGL0X1l
GFzL3xM6feIPRTmW7kgaOCqgMibHBBv10ti9PWXraBg2kP9eHRi7kwiRfW1BoIP2dDTZA+qeban/
INE8EFkx0QEn6Xe3lPjbYwKrfM7ySwTPdIc8cjTOxKtOP0/WaH7MAIeOo7In4igiibbJER1CGarS
AiB4ea41VeNV4vKXUarJRhzTN7gT+0r0Qe/BPazNUliaPJlaKHuXQ/4CG1iNV2pgmjEo9QV9IehY
i2gYgCSShNRLMI2cU12QXqbUlHNmMzK/a/A2eMDicVGfi+1y+KwXmRL03y2eVl0TzvIlrfrOAgrA
mTxekuaZKw3JXpVEfeoDG2qU2h2nUsngSWrNxHdy4ql1GEfiPop9ByyXA0jp/HFndejYLzsQW342
A85SVp/RcEBD467dInnH16Lgl8HZzQ4wagYk7WuQ7UjYG5rOu9J5loEYNbiZWERkPJEVGEWQVtaA
rfvwS+YQIkROYn0yKjE75w3Iosvpchg5kUwLIHm6Uwn+9aFKw3qDU2mpys3vBVFI8sWBGRI0KvGC
oyRcAaNxi3r6wySd8wmjd/UXlqWTlxFMVBwwD5aLd9BjlFk5nzimmnS63DBBdpkZXR6GhcXJvy+u
76MhU6xtF+kXXQSiBtuuR1dSa5K8v4W8h+X7w8xvnwWdWmTXasf/y8pQlKm7lBr3B8OOoip8frVp
JHBc/7l+CTnfkz7nBxpWcKa0+7vjmgGM58+mRZn+iFvVhSP8jLNIs4t7KCf7zJMWUAm3F5oMY2Sh
Gf4jXYAMrr3NI6i0BzChYiXX0GCI859dDQ0VRvl2PUwYNFlEX0DpX7D1Yd6dAzGPRCnuNhIl+z7g
2GfmFC3do5VggagsqvKqRirkIBQD9V9/eezZiy/wH+kSveXaOL9SFMnuoeUo6zSwRtweHHzhAKB0
0SRK7HLzlRuWPJpgwijDuIYjvU3gG/u9u8FoPANG6lQ7EHh31YqGNho4mrI/mUBpO4HbV7IqU4Ty
3Gzrjg72dSry9QwITlsukzTcpnSTNwVa4csfJohL+TDYNwHMgDK3cuvhoAId1ALD1Q+T1CIOCE1r
0un979FyK0KiJJUlSDke9+HPSWPmlW4Ty8XeGWAqgTyeelByCwrU7PitELiFq3t3n4Mvs7957Kkt
SCwzhHQNpG4x+74ej5AOhK/q728xYqsBznaJvOpCcUKAlKtYkkDPjwbvClqfjZdt+7ASk0RjTnkT
H8ldKo67Pah1uMTvwipm2M+EdcU8J884Rsgg1/HqffZ119u8sUOsf7HB5xgW6ekFJZZKfGOAwKe/
tF7UB+RZqIRwdjPfin6ubbt/r74XOK1G/IWB6UoFChJPLxPct1gVuADbfTJkdwtfrGGDLQUry1nE
K+X3PceBVbOgOtmT2nfu6mSDYsS/Dt9VJMQXgB6BuEgebQi1LG1uzl4bd+bO78rq/J7JsN6V3QT+
7UIPMSkPo0AY5ZNXvxpfBAMWqRy2tShHb14lbDOrXV+4YOR1tnIvBHkoWFzHIK5cej8Ri8qGHhg3
NeW9MndpPV6uicP+CXJcp9HVWsUYfpYMCxZb+VrRmKVlK6miePivR27iHi2e7VsoanFYcrxGd7M+
sRlXFL+XzFqeaO2eqo5aoKvLqJsaQgxjK7ItUi9FIweCjVexC/TQO1HRX0fXDRk1Xc9KDc2+/+Uz
aaFQLKBaxAzxHG/Nx/Qdme4oDkrjuq9RPCES4L1TGYuRzNzqtEDR20tok7n4MdG2UTM+1hfQKQ3r
UEy8Z7eHEz0/3YE84iznG11nqYasMT6E4Id6VautKLZZrGKIIy5eqtilEpo5ccCplLrFz9orMxO+
0MTQG+oUMhAr6mPOVAgrWNqBEPkTfN0bEnsYc/T0SjLnwiFMotwzdf8B0PB9CfXPBdSQLoHjuSpM
JMz/GbQ34vtSqtNEjaiC9wZlLlUsdY7EI031R5kyqMlG3Ml078J1DwtrYbJCibG5WUcFtid+bwsL
Q7um9fIuXt7dvfTVS9cZ8NFj9T8tg08AHimeek3kBdz42Q2LLICNTLlMBLIhsicrCZAlFLwcJibc
8rGABzzJnL9Y9IOyBN02c8w+btowELSEoq9V3eNefkVSOwVxdOLsTIwkyKUX8G3cVEPDCkK3WUU/
4B9ucPNhKp94EGEGSeIJIC1QhwWWMyzISz6uCkParQ9mHMwbzYDfM/pctCpId0I9UgHcxwaw1u32
7KX6ASdVpDA4IPkar9xctLQFTtDh3W56PkmdJZB3B2bzJeaPlDxF7d1cuR/7rAAOIq7vcBVXON7L
A96cslztgD6ZOsp3ZhQkBV35CE+XYshGuYsIVzAW1SgvreoNpdZYPWKlVN9jr+iqpwzT8bNjxIyy
oY3KkoCniW2jOkSvn01/K5ApbMHEfYXJv9pWH2/xzNr6G6In4awcgbofqGKvu7+gpQzYrVAKrZ7x
7HnNaYyH3Y+POIz1oF/nkvhEO70Im28xuvlrFFS1yMj/GIjHm4yKHo8yGo8vkyrMJAu3qYlVlk12
nVwXWnJJhC3xV4FJy4PVIB7Ir83efhoqMy8DtDZlKLH6MIrKu4P8+SgOG5SA6mRaDfRAFiTMR+JV
VcX3opHWAiIS9sU1ABmjlvaiB5W9UhbR1X3CJqavxoSnmItqcn/dR43iHfxttSo8KB9FZs4vC8nv
uF57IgWzwa29BAJQAC6BoWUQBkUBDifH8PDLyZVh7tal3m+fNXDH5UtBh3F9/zcow4Nx0W553Eao
zQ2GD08PfqL1StSGMzt/5G5j+27ZcZOBkDVgif2+D4KL7Yhu+PyQJpD1teWtY0p+PbX2ZTJOeAGF
fZW+rGIEgLsg/A41bZOXNvlzY44S97gzdV7qhrI9K+82T3mputWp2iKNYJuzcahBM3vJUbJxtqNB
q+hAf8dE90bW0pYxwlyhcT4uGIT594aEuzp/HWiLf5tjQeAUXHjUIh6W8wEZ0ux3dK9dqmDQx9ia
ZoBO6CV6pNDhvrJXLG6jKMdZc0SLNJIpfsGdV5JWZPEwIzmXC829jIHIlyrP2gx+S/9XNeUxUvkz
l7IS6VqtHl5uTnPLZtK1cuOwW3FnJDlca9jGqM47ChSJUr2ZgvYR1gEDgVmBElZqv0qoUTJvX+Th
0YDPULVVZGU6JFsvmvG5dVWow2NVoDKtw7PqrCGFJZO9ZvW6Bxvqi4+t/u+7llYFp5mIJIsgWw9j
CyJWjdLCGCERBqcE2nMCu8AcX+TgiY8niSvfYh6V3YvlUymv/2vteRpGcx80Y2HNUcLNguCaGB07
rw/tgVg7DHp34SBG03Q4H8V95oeCyljwasO1ZV+TXFrzN2knDgKeRdCw5cp2OPd2R6ihfPkV9aln
fT/CYQzTM7tM5wSSTfWDgLQ87U2rpg==
`pragma protect end_protected
